magic
tech sky130A
magscale 1 2
timestamp 1623893300
<< obsli1 >>
rect 1104 2159 39807 117521
<< obsm1 >>
rect 106 82272 40000 118244
rect 106 82220 40006 82272
rect 106 65068 40000 82220
rect 106 65016 40006 65068
rect 106 1504 40000 65016
<< metal2 >>
rect 110 119200 166 120800
rect 294 119200 350 120800
rect 570 119200 626 120800
rect 754 119200 810 120800
rect 1030 119200 1086 120800
rect 1214 119200 1270 120800
rect 1490 119200 1546 120800
rect 1674 119200 1730 120800
rect 1950 119200 2006 120800
rect 2134 119200 2190 120800
rect 2410 119200 2466 120800
rect 2594 119200 2650 120800
rect 2870 119200 2926 120800
rect 3054 119200 3110 120800
rect 3330 119200 3386 120800
rect 3514 119200 3570 120800
rect 3790 119200 3846 120800
rect 3974 119200 4030 120800
rect 4250 119200 4306 120800
rect 4434 119200 4490 120800
rect 4710 119200 4766 120800
rect 4894 119200 4950 120800
rect 5170 119200 5226 120800
rect 5354 119200 5410 120800
rect 5630 119200 5686 120800
rect 5814 119200 5870 120800
rect 6090 119200 6146 120800
rect 6274 119200 6330 120800
rect 6550 119200 6606 120800
rect 6734 119200 6790 120800
rect 7010 119200 7066 120800
rect 7194 119200 7250 120800
rect 7470 119200 7526 120800
rect 7654 119200 7710 120800
rect 7930 119200 7986 120800
rect 8206 119200 8262 120800
rect 8390 119200 8446 120800
rect 8666 119200 8722 120800
rect 8850 119200 8906 120800
rect 9126 119200 9182 120800
rect 9310 119200 9366 120800
rect 9586 119200 9642 120800
rect 9770 119200 9826 120800
rect 10046 119200 10102 120800
rect 10230 119200 10286 120800
rect 10506 119200 10562 120800
rect 10690 119200 10746 120800
rect 10966 119200 11022 120800
rect 11150 119200 11206 120800
rect 11426 119200 11482 120800
rect 11610 119200 11666 120800
rect 11886 119200 11942 120800
rect 12070 119200 12126 120800
rect 12346 119200 12402 120800
rect 12530 119200 12586 120800
rect 12806 119200 12862 120800
rect 12990 119200 13046 120800
rect 13266 119200 13322 120800
rect 13450 119200 13506 120800
rect 13726 119200 13782 120800
rect 13910 119200 13966 120800
rect 14186 119200 14242 120800
rect 14370 119200 14426 120800
rect 14646 119200 14702 120800
rect 14830 119200 14886 120800
rect 15106 119200 15162 120800
rect 15290 119200 15346 120800
rect 15566 119200 15622 120800
rect 15750 119200 15806 120800
rect 16026 119200 16082 120800
rect 16302 119200 16358 120800
rect 16486 119200 16542 120800
rect 16762 119200 16818 120800
rect 16946 119200 17002 120800
rect 17222 119200 17278 120800
rect 17406 119200 17462 120800
rect 17682 119200 17738 120800
rect 17866 119200 17922 120800
rect 18142 119200 18198 120800
rect 18326 119200 18382 120800
rect 18602 119200 18658 120800
rect 18786 119200 18842 120800
rect 19062 119200 19118 120800
rect 19246 119200 19302 120800
rect 19522 119200 19578 120800
rect 19706 119200 19762 120800
rect 19982 119200 20038 120800
rect 20166 119200 20222 120800
rect 20442 119200 20498 120800
rect 20626 119200 20682 120800
rect 20902 119200 20958 120800
rect 21086 119200 21142 120800
rect 21362 119200 21418 120800
rect 21546 119200 21602 120800
rect 21822 119200 21878 120800
rect 22006 119200 22062 120800
rect 22282 119200 22338 120800
rect 22466 119200 22522 120800
rect 22742 119200 22798 120800
rect 22926 119200 22982 120800
rect 23202 119200 23258 120800
rect 23386 119200 23442 120800
rect 23662 119200 23718 120800
rect 23846 119200 23902 120800
rect 24122 119200 24178 120800
rect 24398 119200 24454 120800
rect 24582 119200 24638 120800
rect 24858 119200 24914 120800
rect 25042 119200 25098 120800
rect 25318 119200 25374 120800
rect 25502 119200 25558 120800
rect 25778 119200 25834 120800
rect 25962 119200 26018 120800
rect 26238 119200 26294 120800
rect 26422 119200 26478 120800
rect 26698 119200 26754 120800
rect 26882 119200 26938 120800
rect 27158 119200 27214 120800
rect 27342 119200 27398 120800
rect 27618 119200 27674 120800
rect 27802 119200 27858 120800
rect 28078 119200 28134 120800
rect 28262 119200 28318 120800
rect 28538 119200 28594 120800
rect 28722 119200 28778 120800
rect 28998 119200 29054 120800
rect 29182 119200 29238 120800
rect 29458 119200 29514 120800
rect 29642 119200 29698 120800
rect 29918 119200 29974 120800
rect 30102 119200 30158 120800
rect 30378 119200 30434 120800
rect 30562 119200 30618 120800
rect 30838 119200 30894 120800
rect 31022 119200 31078 120800
rect 31298 119200 31354 120800
rect 31482 119200 31538 120800
rect 31758 119200 31814 120800
rect 31942 119200 31998 120800
rect 32218 119200 32274 120800
rect 32494 119200 32550 120800
rect 32678 119200 32734 120800
rect 32954 119200 33010 120800
rect 33138 119200 33194 120800
rect 33414 119200 33470 120800
rect 33598 119200 33654 120800
rect 33874 119200 33930 120800
rect 34058 119200 34114 120800
rect 34334 119200 34390 120800
rect 34518 119200 34574 120800
rect 34794 119200 34850 120800
rect 34978 119200 35034 120800
rect 35254 119200 35310 120800
rect 35438 119200 35494 120800
rect 35714 119200 35770 120800
rect 35898 119200 35954 120800
rect 36174 119200 36230 120800
rect 36358 119200 36414 120800
rect 36634 119200 36690 120800
rect 36818 119200 36874 120800
rect 37094 119200 37150 120800
rect 37278 119200 37334 120800
rect 37554 119200 37610 120800
rect 37738 119200 37794 120800
rect 38014 119200 38070 120800
rect 38198 119200 38254 120800
rect 38474 119200 38530 120800
rect 38658 119200 38714 120800
rect 38934 119200 38990 120800
rect 39118 119200 39174 120800
rect 39394 119200 39450 120800
rect 39578 119200 39634 120800
rect 39854 119200 39910 120800
rect 110 -800 166 800
rect 386 -800 442 800
rect 754 -800 810 800
rect 1030 -800 1086 800
rect 1398 -800 1454 800
rect 1674 -800 1730 800
rect 2042 -800 2098 800
rect 2318 -800 2374 800
rect 2686 -800 2742 800
rect 2962 -800 3018 800
rect 3330 -800 3386 800
rect 3606 -800 3662 800
rect 3974 -800 4030 800
rect 4250 -800 4306 800
rect 4618 -800 4674 800
rect 4986 -800 5042 800
rect 5262 -800 5318 800
rect 5630 -800 5686 800
rect 5906 -800 5962 800
rect 6274 -800 6330 800
rect 6550 -800 6606 800
rect 6918 -800 6974 800
rect 7194 -800 7250 800
rect 7562 -800 7618 800
rect 7838 -800 7894 800
rect 8206 -800 8262 800
rect 8482 -800 8538 800
rect 8850 -800 8906 800
rect 9218 -800 9274 800
rect 9494 -800 9550 800
rect 9862 -800 9918 800
rect 10138 -800 10194 800
rect 10506 -800 10562 800
rect 10782 -800 10838 800
rect 11150 -800 11206 800
rect 11426 -800 11482 800
rect 11794 -800 11850 800
rect 12070 -800 12126 800
rect 12438 -800 12494 800
rect 12714 -800 12770 800
rect 13082 -800 13138 800
rect 13450 -800 13506 800
rect 13726 -800 13782 800
rect 14094 -800 14150 800
rect 14370 -800 14426 800
rect 14738 -800 14794 800
rect 15014 -800 15070 800
rect 15382 -800 15438 800
rect 15658 -800 15714 800
rect 16026 -800 16082 800
rect 16302 -800 16358 800
rect 16670 -800 16726 800
rect 16946 -800 17002 800
rect 17314 -800 17370 800
rect 17590 -800 17646 800
rect 17958 -800 18014 800
rect 18326 -800 18382 800
rect 18602 -800 18658 800
rect 18970 -800 19026 800
rect 19246 -800 19302 800
rect 19614 -800 19670 800
rect 19890 -800 19946 800
rect 20258 -800 20314 800
rect 20534 -800 20590 800
rect 20902 -800 20958 800
rect 21178 -800 21234 800
rect 21546 -800 21602 800
rect 21822 -800 21878 800
rect 22190 -800 22246 800
rect 22558 -800 22614 800
rect 22834 -800 22890 800
rect 23202 -800 23258 800
rect 23478 -800 23534 800
rect 23846 -800 23902 800
rect 24122 -800 24178 800
rect 24490 -800 24546 800
rect 24766 -800 24822 800
rect 25134 -800 25190 800
rect 25410 -800 25466 800
rect 25778 -800 25834 800
rect 26054 -800 26110 800
rect 26422 -800 26478 800
rect 26790 -800 26846 800
rect 27066 -800 27122 800
rect 27434 -800 27490 800
rect 27710 -800 27766 800
rect 28078 -800 28134 800
rect 28354 -800 28410 800
rect 28722 -800 28778 800
rect 28998 -800 29054 800
rect 29366 -800 29422 800
rect 29642 -800 29698 800
rect 30010 -800 30066 800
rect 30286 -800 30342 800
rect 30654 -800 30710 800
rect 30930 -800 30986 800
rect 31298 -800 31354 800
rect 31666 -800 31722 800
rect 31942 -800 31998 800
rect 32310 -800 32366 800
rect 32586 -800 32642 800
rect 32954 -800 33010 800
rect 33230 -800 33286 800
rect 33598 -800 33654 800
rect 33874 -800 33930 800
rect 34242 -800 34298 800
rect 34518 -800 34574 800
rect 34886 -800 34942 800
rect 35162 -800 35218 800
rect 35530 -800 35586 800
rect 35898 -800 35954 800
rect 36174 -800 36230 800
rect 36542 -800 36598 800
rect 36818 -800 36874 800
rect 37186 -800 37242 800
rect 37462 -800 37518 800
rect 37830 -800 37886 800
rect 38106 -800 38162 800
rect 38474 -800 38530 800
rect 38750 -800 38806 800
rect 39118 -800 39174 800
rect 39394 -800 39450 800
rect 39762 -800 39818 800
<< obsm2 >>
rect 222 119144 238 119649
rect 406 119144 514 119649
rect 682 119144 698 119649
rect 866 119144 974 119649
rect 1142 119144 1158 119649
rect 1326 119144 1434 119649
rect 1602 119144 1618 119649
rect 1786 119144 1894 119649
rect 2062 119144 2078 119649
rect 2246 119144 2354 119649
rect 2522 119144 2538 119649
rect 2706 119144 2814 119649
rect 2982 119144 2998 119649
rect 3166 119144 3274 119649
rect 3442 119144 3458 119649
rect 3626 119144 3734 119649
rect 3902 119144 3918 119649
rect 4086 119144 4194 119649
rect 4362 119144 4378 119649
rect 4546 119144 4654 119649
rect 4822 119144 4838 119649
rect 5006 119144 5114 119649
rect 5282 119144 5298 119649
rect 5466 119144 5574 119649
rect 5742 119144 5758 119649
rect 5926 119144 6034 119649
rect 6202 119144 6218 119649
rect 6386 119144 6494 119649
rect 6662 119144 6678 119649
rect 6846 119144 6954 119649
rect 7122 119144 7138 119649
rect 7306 119144 7414 119649
rect 7582 119144 7598 119649
rect 7766 119144 7874 119649
rect 8042 119144 8150 119649
rect 8318 119144 8334 119649
rect 8502 119144 8610 119649
rect 8778 119144 8794 119649
rect 8962 119144 9070 119649
rect 9238 119144 9254 119649
rect 9422 119144 9530 119649
rect 9698 119144 9714 119649
rect 9882 119144 9990 119649
rect 10158 119144 10174 119649
rect 10342 119144 10450 119649
rect 10618 119144 10634 119649
rect 10802 119144 10910 119649
rect 11078 119144 11094 119649
rect 11262 119144 11370 119649
rect 11538 119144 11554 119649
rect 11722 119144 11830 119649
rect 11998 119144 12014 119649
rect 12182 119144 12290 119649
rect 12458 119144 12474 119649
rect 12642 119144 12750 119649
rect 12918 119144 12934 119649
rect 13102 119144 13210 119649
rect 13378 119144 13394 119649
rect 13562 119144 13670 119649
rect 13838 119144 13854 119649
rect 14022 119144 14130 119649
rect 14298 119144 14314 119649
rect 14482 119144 14590 119649
rect 14758 119144 14774 119649
rect 14942 119144 15050 119649
rect 15218 119144 15234 119649
rect 15402 119144 15510 119649
rect 15678 119144 15694 119649
rect 15862 119144 15970 119649
rect 16138 119144 16246 119649
rect 16414 119144 16430 119649
rect 16598 119144 16706 119649
rect 16874 119144 16890 119649
rect 17058 119144 17166 119649
rect 17334 119144 17350 119649
rect 17518 119144 17626 119649
rect 17794 119144 17810 119649
rect 17978 119144 18086 119649
rect 18254 119144 18270 119649
rect 18438 119144 18546 119649
rect 18714 119144 18730 119649
rect 18898 119144 19006 119649
rect 19174 119144 19190 119649
rect 19358 119144 19466 119649
rect 19634 119144 19650 119649
rect 19818 119144 19926 119649
rect 20094 119144 20110 119649
rect 20278 119144 20386 119649
rect 20554 119144 20570 119649
rect 20738 119144 20846 119649
rect 21014 119144 21030 119649
rect 21198 119144 21306 119649
rect 21474 119144 21490 119649
rect 21658 119144 21766 119649
rect 21934 119144 21950 119649
rect 22118 119144 22226 119649
rect 22394 119144 22410 119649
rect 22578 119144 22686 119649
rect 22854 119144 22870 119649
rect 23038 119144 23146 119649
rect 23314 119144 23330 119649
rect 23498 119144 23606 119649
rect 23774 119144 23790 119649
rect 23958 119144 24066 119649
rect 24234 119144 24342 119649
rect 24510 119144 24526 119649
rect 24694 119144 24802 119649
rect 24970 119144 24986 119649
rect 25154 119144 25262 119649
rect 25430 119144 25446 119649
rect 25614 119144 25722 119649
rect 25890 119144 25906 119649
rect 26074 119144 26182 119649
rect 26350 119144 26366 119649
rect 26534 119144 26642 119649
rect 26810 119144 26826 119649
rect 26994 119144 27102 119649
rect 27270 119144 27286 119649
rect 27454 119144 27562 119649
rect 27730 119144 27746 119649
rect 27914 119144 28022 119649
rect 28190 119144 28206 119649
rect 28374 119144 28482 119649
rect 28650 119144 28666 119649
rect 28834 119144 28942 119649
rect 29110 119144 29126 119649
rect 29294 119144 29402 119649
rect 29570 119144 29586 119649
rect 29754 119144 29862 119649
rect 30030 119144 30046 119649
rect 30214 119144 30322 119649
rect 30490 119144 30506 119649
rect 30674 119144 30782 119649
rect 30950 119144 30966 119649
rect 31134 119144 31242 119649
rect 31410 119144 31426 119649
rect 31594 119144 31702 119649
rect 31870 119144 31886 119649
rect 32054 119144 32162 119649
rect 32330 119144 32438 119649
rect 32606 119144 32622 119649
rect 32790 119144 32898 119649
rect 33066 119144 33082 119649
rect 33250 119144 33358 119649
rect 33526 119144 33542 119649
rect 33710 119144 33818 119649
rect 33986 119144 34002 119649
rect 34170 119144 34278 119649
rect 34446 119144 34462 119649
rect 34630 119144 34738 119649
rect 34906 119144 34922 119649
rect 35090 119144 35198 119649
rect 35366 119144 35382 119649
rect 35550 119144 35658 119649
rect 35826 119144 35842 119649
rect 36010 119144 36118 119649
rect 36286 119144 36302 119649
rect 36470 119144 36578 119649
rect 36746 119144 36762 119649
rect 36930 119144 37038 119649
rect 37206 119144 37222 119649
rect 37390 119144 37498 119649
rect 37666 119144 37682 119649
rect 37850 119144 37958 119649
rect 38126 119144 38142 119649
rect 38310 119144 38418 119649
rect 38586 119144 38602 119649
rect 38770 119144 38878 119649
rect 39046 119144 39062 119649
rect 39230 119144 39338 119649
rect 39506 119144 39522 119649
rect 39690 119144 39798 119649
rect 39966 119144 40000 119649
rect 112 856 40000 119144
rect 222 167 330 856
rect 498 167 698 856
rect 866 167 974 856
rect 1142 167 1342 856
rect 1510 167 1618 856
rect 1786 167 1986 856
rect 2154 167 2262 856
rect 2430 167 2630 856
rect 2798 167 2906 856
rect 3074 167 3274 856
rect 3442 167 3550 856
rect 3718 167 3918 856
rect 4086 167 4194 856
rect 4362 167 4562 856
rect 4730 167 4930 856
rect 5098 167 5206 856
rect 5374 167 5574 856
rect 5742 167 5850 856
rect 6018 167 6218 856
rect 6386 167 6494 856
rect 6662 167 6862 856
rect 7030 167 7138 856
rect 7306 167 7506 856
rect 7674 167 7782 856
rect 7950 167 8150 856
rect 8318 167 8426 856
rect 8594 167 8794 856
rect 8962 167 9162 856
rect 9330 167 9438 856
rect 9606 167 9806 856
rect 9974 167 10082 856
rect 10250 167 10450 856
rect 10618 167 10726 856
rect 10894 167 11094 856
rect 11262 167 11370 856
rect 11538 167 11738 856
rect 11906 167 12014 856
rect 12182 167 12382 856
rect 12550 167 12658 856
rect 12826 167 13026 856
rect 13194 167 13394 856
rect 13562 167 13670 856
rect 13838 167 14038 856
rect 14206 167 14314 856
rect 14482 167 14682 856
rect 14850 167 14958 856
rect 15126 167 15326 856
rect 15494 167 15602 856
rect 15770 167 15970 856
rect 16138 167 16246 856
rect 16414 167 16614 856
rect 16782 167 16890 856
rect 17058 167 17258 856
rect 17426 167 17534 856
rect 17702 167 17902 856
rect 18070 167 18270 856
rect 18438 167 18546 856
rect 18714 167 18914 856
rect 19082 167 19190 856
rect 19358 167 19558 856
rect 19726 167 19834 856
rect 20002 167 20202 856
rect 20370 167 20478 856
rect 20646 167 20846 856
rect 21014 167 21122 856
rect 21290 167 21490 856
rect 21658 167 21766 856
rect 21934 167 22134 856
rect 22302 167 22502 856
rect 22670 167 22778 856
rect 22946 167 23146 856
rect 23314 167 23422 856
rect 23590 167 23790 856
rect 23958 167 24066 856
rect 24234 167 24434 856
rect 24602 167 24710 856
rect 24878 167 25078 856
rect 25246 167 25354 856
rect 25522 167 25722 856
rect 25890 167 25998 856
rect 26166 167 26366 856
rect 26534 167 26734 856
rect 26902 167 27010 856
rect 27178 167 27378 856
rect 27546 167 27654 856
rect 27822 167 28022 856
rect 28190 167 28298 856
rect 28466 167 28666 856
rect 28834 167 28942 856
rect 29110 167 29310 856
rect 29478 167 29586 856
rect 29754 167 29954 856
rect 30122 167 30230 856
rect 30398 167 30598 856
rect 30766 167 30874 856
rect 31042 167 31242 856
rect 31410 167 31610 856
rect 31778 167 31886 856
rect 32054 167 32254 856
rect 32422 167 32530 856
rect 32698 167 32898 856
rect 33066 167 33174 856
rect 33342 167 33542 856
rect 33710 167 33818 856
rect 33986 167 34186 856
rect 34354 167 34462 856
rect 34630 167 34830 856
rect 34998 167 35106 856
rect 35274 167 35474 856
rect 35642 167 35842 856
rect 36010 167 36118 856
rect 36286 167 36486 856
rect 36654 167 36762 856
rect 36930 167 37130 856
rect 37298 167 37406 856
rect 37574 167 37774 856
rect 37942 167 38050 856
rect 38218 167 38418 856
rect 38586 167 38694 856
rect 38862 167 39062 856
rect 39230 167 39338 856
rect 39506 167 39706 856
rect 39874 167 40000 856
<< metal3 >>
rect -800 119416 800 119536
rect 39200 119552 40800 119672
rect 39200 119144 40800 119264
rect -800 118600 800 118720
rect 39200 118736 40800 118856
rect 39200 118192 40800 118312
rect -800 117784 800 117904
rect 39200 117784 40800 117904
rect 39200 117376 40800 117496
rect -800 116968 800 117088
rect 39200 116832 40800 116952
rect 39200 116424 40800 116544
rect -800 116152 800 116272
rect 39200 116016 40800 116136
rect 39200 115608 40800 115728
rect -800 115336 800 115456
rect 39200 115064 40800 115184
rect -800 114520 800 114640
rect 39200 114656 40800 114776
rect 39200 114248 40800 114368
rect -800 113704 800 113824
rect 39200 113704 40800 113824
rect 39200 113296 40800 113416
rect -800 113024 800 113144
rect 39200 112888 40800 113008
rect 39200 112480 40800 112600
rect -800 112208 800 112328
rect 39200 111936 40800 112056
rect -800 111392 800 111512
rect 39200 111528 40800 111648
rect 39200 111120 40800 111240
rect -800 110576 800 110696
rect 39200 110576 40800 110696
rect 39200 110168 40800 110288
rect -800 109760 800 109880
rect 39200 109760 40800 109880
rect 39200 109352 40800 109472
rect -800 108944 800 109064
rect 39200 108808 40800 108928
rect 39200 108400 40800 108520
rect -800 108128 800 108248
rect 39200 107992 40800 108112
rect -800 107312 800 107432
rect 39200 107448 40800 107568
rect 39200 107040 40800 107160
rect -800 106632 800 106752
rect 39200 106632 40800 106752
rect 39200 106088 40800 106208
rect -800 105816 800 105936
rect 39200 105680 40800 105800
rect 39200 105272 40800 105392
rect -800 105000 800 105120
rect 39200 104864 40800 104984
rect -800 104184 800 104304
rect 39200 104320 40800 104440
rect 39200 103912 40800 104032
rect -800 103368 800 103488
rect 39200 103504 40800 103624
rect 39200 102960 40800 103080
rect -800 102552 800 102672
rect 39200 102552 40800 102672
rect 39200 102144 40800 102264
rect -800 101736 800 101856
rect 39200 101736 40800 101856
rect 39200 101192 40800 101312
rect -800 100920 800 101040
rect 39200 100784 40800 100904
rect -800 100240 800 100360
rect 39200 100376 40800 100496
rect 39200 99832 40800 99952
rect -800 99424 800 99544
rect 39200 99424 40800 99544
rect 39200 99016 40800 99136
rect -800 98608 800 98728
rect 39200 98608 40800 98728
rect 39200 98064 40800 98184
rect -800 97792 800 97912
rect 39200 97656 40800 97776
rect 39200 97248 40800 97368
rect -800 96976 800 97096
rect 39200 96704 40800 96824
rect -800 96160 800 96280
rect 39200 96296 40800 96416
rect 39200 95888 40800 96008
rect -800 95344 800 95464
rect 39200 95344 40800 95464
rect 39200 94936 40800 95056
rect -800 94528 800 94648
rect 39200 94528 40800 94648
rect 39200 94120 40800 94240
rect -800 93712 800 93832
rect 39200 93576 40800 93696
rect -800 93032 800 93152
rect 39200 93168 40800 93288
rect 39200 92760 40800 92880
rect -800 92216 800 92336
rect 39200 92216 40800 92336
rect 39200 91808 40800 91928
rect -800 91400 800 91520
rect 39200 91400 40800 91520
rect 39200 90992 40800 91112
rect -800 90584 800 90704
rect 39200 90448 40800 90568
rect 39200 90040 40800 90160
rect -800 89768 800 89888
rect 39200 89632 40800 89752
rect -800 88952 800 89072
rect 39200 89088 40800 89208
rect 39200 88680 40800 88800
rect -800 88136 800 88256
rect 39200 88272 40800 88392
rect 39200 87864 40800 87984
rect -800 87320 800 87440
rect 39200 87320 40800 87440
rect 39200 86912 40800 87032
rect -800 86640 800 86760
rect 39200 86504 40800 86624
rect -800 85824 800 85944
rect 39200 85960 40800 86080
rect 39200 85552 40800 85672
rect -800 85008 800 85128
rect 39200 85144 40800 85264
rect 39200 84736 40800 84856
rect -800 84192 800 84312
rect 39200 84192 40800 84312
rect 39200 83784 40800 83904
rect -800 83376 800 83496
rect 39200 83376 40800 83496
rect 39200 82832 40800 82952
rect -800 82560 800 82680
rect 39200 82424 40800 82544
rect 39200 82016 40800 82136
rect -800 81744 800 81864
rect 39200 81472 40800 81592
rect -800 80928 800 81048
rect 39200 81064 40800 81184
rect 39200 80656 40800 80776
rect -800 80248 800 80368
rect 39200 80248 40800 80368
rect 39200 79704 40800 79824
rect -800 79432 800 79552
rect 39200 79296 40800 79416
rect 39200 78888 40800 79008
rect -800 78616 800 78736
rect 39200 78344 40800 78464
rect -800 77800 800 77920
rect 39200 77936 40800 78056
rect 39200 77528 40800 77648
rect -800 76984 800 77104
rect 39200 77120 40800 77240
rect 39200 76576 40800 76696
rect -800 76168 800 76288
rect 39200 76168 40800 76288
rect 39200 75760 40800 75880
rect -800 75352 800 75472
rect 39200 75216 40800 75336
rect 39200 74808 40800 74928
rect -800 74536 800 74656
rect 39200 74400 40800 74520
rect 39200 73992 40800 74112
rect -800 73720 800 73840
rect 39200 73448 40800 73568
rect -800 73040 800 73160
rect 39200 73040 40800 73160
rect 39200 72632 40800 72752
rect -800 72224 800 72344
rect 39200 72088 40800 72208
rect 39200 71680 40800 71800
rect -800 71408 800 71528
rect 39200 71272 40800 71392
rect -800 70592 800 70712
rect 39200 70728 40800 70848
rect 39200 70320 40800 70440
rect -800 69776 800 69896
rect 39200 69912 40800 70032
rect 39200 69504 40800 69624
rect -800 68960 800 69080
rect 39200 68960 40800 69080
rect 39200 68552 40800 68672
rect -800 68144 800 68264
rect 39200 68144 40800 68264
rect 39200 67600 40800 67720
rect -800 67328 800 67448
rect 39200 67192 40800 67312
rect -800 66648 800 66768
rect 39200 66784 40800 66904
rect 39200 66376 40800 66496
rect -800 65832 800 65952
rect 39200 65832 40800 65952
rect 39200 65424 40800 65544
rect -800 65016 800 65136
rect 39200 65016 40800 65136
rect 39200 64472 40800 64592
rect -800 64200 800 64320
rect 39200 64064 40800 64184
rect 39200 63656 40800 63776
rect -800 63384 800 63504
rect 39200 63248 40800 63368
rect -800 62568 800 62688
rect 39200 62704 40800 62824
rect 39200 62296 40800 62416
rect -800 61752 800 61872
rect 39200 61888 40800 62008
rect 39200 61344 40800 61464
rect -800 60936 800 61056
rect 39200 60936 40800 61056
rect 39200 60528 40800 60648
rect -800 60256 800 60376
rect 39200 60120 40800 60240
rect -800 59440 800 59560
rect 39200 59576 40800 59696
rect 39200 59168 40800 59288
rect -800 58624 800 58744
rect 39200 58760 40800 58880
rect 39200 58216 40800 58336
rect -800 57808 800 57928
rect 39200 57808 40800 57928
rect 39200 57400 40800 57520
rect -800 56992 800 57112
rect 39200 56856 40800 56976
rect 39200 56448 40800 56568
rect -800 56176 800 56296
rect 39200 56040 40800 56160
rect 39200 55632 40800 55752
rect -800 55360 800 55480
rect 39200 55088 40800 55208
rect -800 54544 800 54664
rect 39200 54680 40800 54800
rect 39200 54272 40800 54392
rect -800 53728 800 53848
rect 39200 53728 40800 53848
rect 39200 53320 40800 53440
rect -800 53048 800 53168
rect 39200 52912 40800 53032
rect 39200 52504 40800 52624
rect -800 52232 800 52352
rect 39200 51960 40800 52080
rect -800 51416 800 51536
rect 39200 51552 40800 51672
rect 39200 51144 40800 51264
rect -800 50600 800 50720
rect 39200 50600 40800 50720
rect 39200 50192 40800 50312
rect -800 49784 800 49904
rect 39200 49784 40800 49904
rect 39200 49376 40800 49496
rect -800 48968 800 49088
rect 39200 48832 40800 48952
rect 39200 48424 40800 48544
rect -800 48152 800 48272
rect 39200 48016 40800 48136
rect -800 47336 800 47456
rect 39200 47472 40800 47592
rect 39200 47064 40800 47184
rect -800 46656 800 46776
rect 39200 46656 40800 46776
rect 39200 46112 40800 46232
rect -800 45840 800 45960
rect 39200 45704 40800 45824
rect 39200 45296 40800 45416
rect -800 45024 800 45144
rect 39200 44888 40800 45008
rect -800 44208 800 44328
rect 39200 44344 40800 44464
rect 39200 43936 40800 44056
rect -800 43392 800 43512
rect 39200 43528 40800 43648
rect 39200 42984 40800 43104
rect -800 42576 800 42696
rect 39200 42576 40800 42696
rect 39200 42168 40800 42288
rect -800 41760 800 41880
rect 39200 41760 40800 41880
rect 39200 41216 40800 41336
rect -800 40944 800 41064
rect 39200 40808 40800 40928
rect -800 40264 800 40384
rect 39200 40400 40800 40520
rect 39200 39856 40800 39976
rect -800 39448 800 39568
rect 39200 39448 40800 39568
rect 39200 39040 40800 39160
rect -800 38632 800 38752
rect 39200 38632 40800 38752
rect 39200 38088 40800 38208
rect -800 37816 800 37936
rect 39200 37680 40800 37800
rect 39200 37272 40800 37392
rect -800 37000 800 37120
rect 39200 36728 40800 36848
rect -800 36184 800 36304
rect 39200 36320 40800 36440
rect 39200 35912 40800 36032
rect -800 35368 800 35488
rect 39200 35368 40800 35488
rect 39200 34960 40800 35080
rect -800 34552 800 34672
rect 39200 34552 40800 34672
rect 39200 34144 40800 34264
rect -800 33736 800 33856
rect 39200 33600 40800 33720
rect -800 33056 800 33176
rect 39200 33192 40800 33312
rect 39200 32784 40800 32904
rect -800 32240 800 32360
rect 39200 32240 40800 32360
rect 39200 31832 40800 31952
rect -800 31424 800 31544
rect 39200 31424 40800 31544
rect 39200 31016 40800 31136
rect -800 30608 800 30728
rect 39200 30472 40800 30592
rect 39200 30064 40800 30184
rect -800 29792 800 29912
rect 39200 29656 40800 29776
rect -800 28976 800 29096
rect 39200 29112 40800 29232
rect 39200 28704 40800 28824
rect -800 28160 800 28280
rect 39200 28296 40800 28416
rect 39200 27888 40800 28008
rect -800 27344 800 27464
rect 39200 27344 40800 27464
rect 39200 26936 40800 27056
rect -800 26664 800 26784
rect 39200 26528 40800 26648
rect -800 25848 800 25968
rect 39200 25984 40800 26104
rect 39200 25576 40800 25696
rect -800 25032 800 25152
rect 39200 25168 40800 25288
rect 39200 24760 40800 24880
rect -800 24216 800 24336
rect 39200 24216 40800 24336
rect 39200 23808 40800 23928
rect -800 23400 800 23520
rect 39200 23400 40800 23520
rect 39200 22856 40800 22976
rect -800 22584 800 22704
rect 39200 22448 40800 22568
rect 39200 22040 40800 22160
rect -800 21768 800 21888
rect 39200 21496 40800 21616
rect -800 20952 800 21072
rect 39200 21088 40800 21208
rect 39200 20680 40800 20800
rect -800 20272 800 20392
rect 39200 20272 40800 20392
rect 39200 19728 40800 19848
rect -800 19456 800 19576
rect 39200 19320 40800 19440
rect 39200 18912 40800 19032
rect -800 18640 800 18760
rect 39200 18368 40800 18488
rect -800 17824 800 17944
rect 39200 17960 40800 18080
rect 39200 17552 40800 17672
rect -800 17008 800 17128
rect 39200 17144 40800 17264
rect 39200 16600 40800 16720
rect -800 16192 800 16312
rect 39200 16192 40800 16312
rect 39200 15784 40800 15904
rect -800 15376 800 15496
rect 39200 15240 40800 15360
rect 39200 14832 40800 14952
rect -800 14560 800 14680
rect 39200 14424 40800 14544
rect 39200 14016 40800 14136
rect -800 13744 800 13864
rect 39200 13472 40800 13592
rect -800 13064 800 13184
rect 39200 13064 40800 13184
rect 39200 12656 40800 12776
rect -800 12248 800 12368
rect 39200 12112 40800 12232
rect 39200 11704 40800 11824
rect -800 11432 800 11552
rect 39200 11296 40800 11416
rect -800 10616 800 10736
rect 39200 10752 40800 10872
rect 39200 10344 40800 10464
rect -800 9800 800 9920
rect 39200 9936 40800 10056
rect 39200 9528 40800 9648
rect -800 8984 800 9104
rect 39200 8984 40800 9104
rect 39200 8576 40800 8696
rect -800 8168 800 8288
rect 39200 8168 40800 8288
rect 39200 7624 40800 7744
rect -800 7352 800 7472
rect 39200 7216 40800 7336
rect -800 6672 800 6792
rect 39200 6808 40800 6928
rect 39200 6400 40800 6520
rect -800 5856 800 5976
rect 39200 5856 40800 5976
rect 39200 5448 40800 5568
rect -800 5040 800 5160
rect 39200 5040 40800 5160
rect 39200 4496 40800 4616
rect -800 4224 800 4344
rect 39200 4088 40800 4208
rect 39200 3680 40800 3800
rect -800 3408 800 3528
rect 39200 3272 40800 3392
rect -800 2592 800 2712
rect 39200 2728 40800 2848
rect 39200 2320 40800 2440
rect -800 1776 800 1896
rect 39200 1912 40800 2032
rect 39200 1368 40800 1488
rect -800 960 800 1080
rect 39200 960 40800 1080
rect 39200 552 40800 672
rect -800 280 800 400
rect 39200 144 40800 264
<< obsm3 >>
rect 800 119616 39120 119645
rect 880 119472 39120 119616
rect 880 119344 39823 119472
rect 880 119336 39120 119344
rect 800 119064 39120 119336
rect 800 118936 39823 119064
rect 800 118800 39120 118936
rect 880 118656 39120 118800
rect 880 118520 39823 118656
rect 800 118392 39823 118520
rect 800 118112 39120 118392
rect 800 117984 39823 118112
rect 880 117704 39120 117984
rect 800 117576 39823 117704
rect 800 117296 39120 117576
rect 800 117168 39823 117296
rect 880 117032 39823 117168
rect 880 116888 39120 117032
rect 800 116752 39120 116888
rect 800 116624 39823 116752
rect 800 116352 39120 116624
rect 880 116344 39120 116352
rect 880 116216 39823 116344
rect 880 116072 39120 116216
rect 800 115936 39120 116072
rect 800 115808 39823 115936
rect 800 115536 39120 115808
rect 880 115528 39120 115536
rect 880 115264 39823 115528
rect 880 115256 39120 115264
rect 800 114984 39120 115256
rect 800 114856 39823 114984
rect 800 114720 39120 114856
rect 880 114576 39120 114720
rect 880 114448 39823 114576
rect 880 114440 39120 114448
rect 800 114168 39120 114440
rect 800 113904 39823 114168
rect 880 113624 39120 113904
rect 800 113496 39823 113624
rect 800 113224 39120 113496
rect 880 113216 39120 113224
rect 880 113088 39823 113216
rect 880 112944 39120 113088
rect 800 112808 39120 112944
rect 800 112680 39823 112808
rect 800 112408 39120 112680
rect 880 112400 39120 112408
rect 880 112136 39823 112400
rect 880 112128 39120 112136
rect 800 111856 39120 112128
rect 800 111728 39823 111856
rect 800 111592 39120 111728
rect 880 111448 39120 111592
rect 880 111320 39823 111448
rect 880 111312 39120 111320
rect 800 111040 39120 111312
rect 800 110776 39823 111040
rect 880 110496 39120 110776
rect 800 110368 39823 110496
rect 800 110088 39120 110368
rect 800 109960 39823 110088
rect 880 109680 39120 109960
rect 800 109552 39823 109680
rect 800 109272 39120 109552
rect 800 109144 39823 109272
rect 880 109008 39823 109144
rect 880 108864 39120 109008
rect 800 108728 39120 108864
rect 800 108600 39823 108728
rect 800 108328 39120 108600
rect 880 108320 39120 108328
rect 880 108192 39823 108320
rect 880 108048 39120 108192
rect 800 107912 39120 108048
rect 800 107648 39823 107912
rect 800 107512 39120 107648
rect 880 107368 39120 107512
rect 880 107240 39823 107368
rect 880 107232 39120 107240
rect 800 106960 39120 107232
rect 800 106832 39823 106960
rect 880 106552 39120 106832
rect 800 106288 39823 106552
rect 800 106016 39120 106288
rect 880 106008 39120 106016
rect 880 105880 39823 106008
rect 880 105736 39120 105880
rect 800 105600 39120 105736
rect 800 105472 39823 105600
rect 800 105200 39120 105472
rect 880 105192 39120 105200
rect 880 105064 39823 105192
rect 880 104920 39120 105064
rect 800 104784 39120 104920
rect 800 104520 39823 104784
rect 800 104384 39120 104520
rect 880 104240 39120 104384
rect 880 104112 39823 104240
rect 880 104104 39120 104112
rect 800 103832 39120 104104
rect 800 103704 39823 103832
rect 800 103568 39120 103704
rect 880 103424 39120 103568
rect 880 103288 39823 103424
rect 800 103160 39823 103288
rect 800 102880 39120 103160
rect 800 102752 39823 102880
rect 880 102472 39120 102752
rect 800 102344 39823 102472
rect 800 102064 39120 102344
rect 800 101936 39823 102064
rect 880 101656 39120 101936
rect 800 101392 39823 101656
rect 800 101120 39120 101392
rect 880 101112 39120 101120
rect 880 100984 39823 101112
rect 880 100840 39120 100984
rect 800 100704 39120 100840
rect 800 100576 39823 100704
rect 800 100440 39120 100576
rect 880 100296 39120 100440
rect 880 100160 39823 100296
rect 800 100032 39823 100160
rect 800 99752 39120 100032
rect 800 99624 39823 99752
rect 880 99344 39120 99624
rect 800 99216 39823 99344
rect 800 98936 39120 99216
rect 800 98808 39823 98936
rect 880 98528 39120 98808
rect 800 98264 39823 98528
rect 800 97992 39120 98264
rect 880 97984 39120 97992
rect 880 97856 39823 97984
rect 880 97712 39120 97856
rect 800 97576 39120 97712
rect 800 97448 39823 97576
rect 800 97176 39120 97448
rect 880 97168 39120 97176
rect 880 96904 39823 97168
rect 880 96896 39120 96904
rect 800 96624 39120 96896
rect 800 96496 39823 96624
rect 800 96360 39120 96496
rect 880 96216 39120 96360
rect 880 96088 39823 96216
rect 880 96080 39120 96088
rect 800 95808 39120 96080
rect 800 95544 39823 95808
rect 880 95264 39120 95544
rect 800 95136 39823 95264
rect 800 94856 39120 95136
rect 800 94728 39823 94856
rect 880 94448 39120 94728
rect 800 94320 39823 94448
rect 800 94040 39120 94320
rect 800 93912 39823 94040
rect 880 93776 39823 93912
rect 880 93632 39120 93776
rect 800 93496 39120 93632
rect 800 93368 39823 93496
rect 800 93232 39120 93368
rect 880 93088 39120 93232
rect 880 92960 39823 93088
rect 880 92952 39120 92960
rect 800 92680 39120 92952
rect 800 92416 39823 92680
rect 880 92136 39120 92416
rect 800 92008 39823 92136
rect 800 91728 39120 92008
rect 800 91600 39823 91728
rect 880 91320 39120 91600
rect 800 91192 39823 91320
rect 800 90912 39120 91192
rect 800 90784 39823 90912
rect 880 90648 39823 90784
rect 880 90504 39120 90648
rect 800 90368 39120 90504
rect 800 90240 39823 90368
rect 800 89968 39120 90240
rect 880 89960 39120 89968
rect 880 89832 39823 89960
rect 880 89688 39120 89832
rect 800 89552 39120 89688
rect 800 89288 39823 89552
rect 800 89152 39120 89288
rect 880 89008 39120 89152
rect 880 88880 39823 89008
rect 880 88872 39120 88880
rect 800 88600 39120 88872
rect 800 88472 39823 88600
rect 800 88336 39120 88472
rect 880 88192 39120 88336
rect 880 88064 39823 88192
rect 880 88056 39120 88064
rect 800 87784 39120 88056
rect 800 87520 39823 87784
rect 880 87240 39120 87520
rect 800 87112 39823 87240
rect 800 86840 39120 87112
rect 880 86832 39120 86840
rect 880 86704 39823 86832
rect 880 86560 39120 86704
rect 800 86424 39120 86560
rect 800 86160 39823 86424
rect 800 86024 39120 86160
rect 880 85880 39120 86024
rect 880 85752 39823 85880
rect 880 85744 39120 85752
rect 800 85472 39120 85744
rect 800 85344 39823 85472
rect 800 85208 39120 85344
rect 880 85064 39120 85208
rect 880 84936 39823 85064
rect 880 84928 39120 84936
rect 800 84656 39120 84928
rect 800 84392 39823 84656
rect 880 84112 39120 84392
rect 800 83984 39823 84112
rect 800 83704 39120 83984
rect 800 83576 39823 83704
rect 880 83296 39120 83576
rect 800 83032 39823 83296
rect 800 82760 39120 83032
rect 880 82752 39120 82760
rect 880 82624 39823 82752
rect 880 82480 39120 82624
rect 800 82344 39120 82480
rect 800 82216 39823 82344
rect 800 81944 39120 82216
rect 880 81936 39120 81944
rect 880 81672 39823 81936
rect 880 81664 39120 81672
rect 800 81392 39120 81664
rect 800 81264 39823 81392
rect 800 81128 39120 81264
rect 880 80984 39120 81128
rect 880 80856 39823 80984
rect 880 80848 39120 80856
rect 800 80576 39120 80848
rect 800 80448 39823 80576
rect 880 80168 39120 80448
rect 800 79904 39823 80168
rect 800 79632 39120 79904
rect 880 79624 39120 79632
rect 880 79496 39823 79624
rect 880 79352 39120 79496
rect 800 79216 39120 79352
rect 800 79088 39823 79216
rect 800 78816 39120 79088
rect 880 78808 39120 78816
rect 880 78544 39823 78808
rect 880 78536 39120 78544
rect 800 78264 39120 78536
rect 800 78136 39823 78264
rect 800 78000 39120 78136
rect 880 77856 39120 78000
rect 880 77728 39823 77856
rect 880 77720 39120 77728
rect 800 77448 39120 77720
rect 800 77320 39823 77448
rect 800 77184 39120 77320
rect 880 77040 39120 77184
rect 880 76904 39823 77040
rect 800 76776 39823 76904
rect 800 76496 39120 76776
rect 800 76368 39823 76496
rect 880 76088 39120 76368
rect 800 75960 39823 76088
rect 800 75680 39120 75960
rect 800 75552 39823 75680
rect 880 75416 39823 75552
rect 880 75272 39120 75416
rect 800 75136 39120 75272
rect 800 75008 39823 75136
rect 800 74736 39120 75008
rect 880 74728 39120 74736
rect 880 74600 39823 74728
rect 880 74456 39120 74600
rect 800 74320 39120 74456
rect 800 74192 39823 74320
rect 800 73920 39120 74192
rect 880 73912 39120 73920
rect 880 73648 39823 73912
rect 880 73640 39120 73648
rect 800 73368 39120 73640
rect 800 73240 39823 73368
rect 880 72960 39120 73240
rect 800 72832 39823 72960
rect 800 72552 39120 72832
rect 800 72424 39823 72552
rect 880 72288 39823 72424
rect 880 72144 39120 72288
rect 800 72008 39120 72144
rect 800 71880 39823 72008
rect 800 71608 39120 71880
rect 880 71600 39120 71608
rect 880 71472 39823 71600
rect 880 71328 39120 71472
rect 800 71192 39120 71328
rect 800 70928 39823 71192
rect 800 70792 39120 70928
rect 880 70648 39120 70792
rect 880 70520 39823 70648
rect 880 70512 39120 70520
rect 800 70240 39120 70512
rect 800 70112 39823 70240
rect 800 69976 39120 70112
rect 880 69832 39120 69976
rect 880 69704 39823 69832
rect 880 69696 39120 69704
rect 800 69424 39120 69696
rect 800 69160 39823 69424
rect 880 68880 39120 69160
rect 800 68752 39823 68880
rect 800 68472 39120 68752
rect 800 68344 39823 68472
rect 880 68064 39120 68344
rect 800 67800 39823 68064
rect 800 67528 39120 67800
rect 880 67520 39120 67528
rect 880 67392 39823 67520
rect 880 67248 39120 67392
rect 800 67112 39120 67248
rect 800 66984 39823 67112
rect 800 66848 39120 66984
rect 880 66704 39120 66848
rect 880 66576 39823 66704
rect 880 66568 39120 66576
rect 800 66296 39120 66568
rect 800 66032 39823 66296
rect 880 65752 39120 66032
rect 800 65624 39823 65752
rect 800 65344 39120 65624
rect 800 65216 39823 65344
rect 880 64936 39120 65216
rect 800 64672 39823 64936
rect 800 64400 39120 64672
rect 880 64392 39120 64400
rect 880 64264 39823 64392
rect 880 64120 39120 64264
rect 800 63984 39120 64120
rect 800 63856 39823 63984
rect 800 63584 39120 63856
rect 880 63576 39120 63584
rect 880 63448 39823 63576
rect 880 63304 39120 63448
rect 800 63168 39120 63304
rect 800 62904 39823 63168
rect 800 62768 39120 62904
rect 880 62624 39120 62768
rect 880 62496 39823 62624
rect 880 62488 39120 62496
rect 800 62216 39120 62488
rect 800 62088 39823 62216
rect 800 61952 39120 62088
rect 880 61808 39120 61952
rect 880 61672 39823 61808
rect 800 61544 39823 61672
rect 800 61264 39120 61544
rect 800 61136 39823 61264
rect 880 60856 39120 61136
rect 800 60728 39823 60856
rect 800 60456 39120 60728
rect 880 60448 39120 60456
rect 880 60320 39823 60448
rect 880 60176 39120 60320
rect 800 60040 39120 60176
rect 800 59776 39823 60040
rect 800 59640 39120 59776
rect 880 59496 39120 59640
rect 880 59368 39823 59496
rect 880 59360 39120 59368
rect 800 59088 39120 59360
rect 800 58960 39823 59088
rect 800 58824 39120 58960
rect 880 58680 39120 58824
rect 880 58544 39823 58680
rect 800 58416 39823 58544
rect 800 58136 39120 58416
rect 800 58008 39823 58136
rect 880 57728 39120 58008
rect 800 57600 39823 57728
rect 800 57320 39120 57600
rect 800 57192 39823 57320
rect 880 57056 39823 57192
rect 880 56912 39120 57056
rect 800 56776 39120 56912
rect 800 56648 39823 56776
rect 800 56376 39120 56648
rect 880 56368 39120 56376
rect 880 56240 39823 56368
rect 880 56096 39120 56240
rect 800 55960 39120 56096
rect 800 55832 39823 55960
rect 800 55560 39120 55832
rect 880 55552 39120 55560
rect 880 55288 39823 55552
rect 880 55280 39120 55288
rect 800 55008 39120 55280
rect 800 54880 39823 55008
rect 800 54744 39120 54880
rect 880 54600 39120 54744
rect 880 54472 39823 54600
rect 880 54464 39120 54472
rect 800 54192 39120 54464
rect 800 53928 39823 54192
rect 880 53648 39120 53928
rect 800 53520 39823 53648
rect 800 53248 39120 53520
rect 880 53240 39120 53248
rect 880 53112 39823 53240
rect 880 52968 39120 53112
rect 800 52832 39120 52968
rect 800 52704 39823 52832
rect 800 52432 39120 52704
rect 880 52424 39120 52432
rect 880 52160 39823 52424
rect 880 52152 39120 52160
rect 800 51880 39120 52152
rect 800 51752 39823 51880
rect 800 51616 39120 51752
rect 880 51472 39120 51616
rect 880 51344 39823 51472
rect 880 51336 39120 51344
rect 800 51064 39120 51336
rect 800 50800 39823 51064
rect 880 50520 39120 50800
rect 800 50392 39823 50520
rect 800 50112 39120 50392
rect 800 49984 39823 50112
rect 880 49704 39120 49984
rect 800 49576 39823 49704
rect 800 49296 39120 49576
rect 800 49168 39823 49296
rect 880 49032 39823 49168
rect 880 48888 39120 49032
rect 800 48752 39120 48888
rect 800 48624 39823 48752
rect 800 48352 39120 48624
rect 880 48344 39120 48352
rect 880 48216 39823 48344
rect 880 48072 39120 48216
rect 800 47936 39120 48072
rect 800 47672 39823 47936
rect 800 47536 39120 47672
rect 880 47392 39120 47536
rect 880 47264 39823 47392
rect 880 47256 39120 47264
rect 800 46984 39120 47256
rect 800 46856 39823 46984
rect 880 46576 39120 46856
rect 800 46312 39823 46576
rect 800 46040 39120 46312
rect 880 46032 39120 46040
rect 880 45904 39823 46032
rect 880 45760 39120 45904
rect 800 45624 39120 45760
rect 800 45496 39823 45624
rect 800 45224 39120 45496
rect 880 45216 39120 45224
rect 880 45088 39823 45216
rect 880 44944 39120 45088
rect 800 44808 39120 44944
rect 800 44544 39823 44808
rect 800 44408 39120 44544
rect 880 44264 39120 44408
rect 880 44136 39823 44264
rect 880 44128 39120 44136
rect 800 43856 39120 44128
rect 800 43728 39823 43856
rect 800 43592 39120 43728
rect 880 43448 39120 43592
rect 880 43312 39823 43448
rect 800 43184 39823 43312
rect 800 42904 39120 43184
rect 800 42776 39823 42904
rect 880 42496 39120 42776
rect 800 42368 39823 42496
rect 800 42088 39120 42368
rect 800 41960 39823 42088
rect 880 41680 39120 41960
rect 800 41416 39823 41680
rect 800 41144 39120 41416
rect 880 41136 39120 41144
rect 880 41008 39823 41136
rect 880 40864 39120 41008
rect 800 40728 39120 40864
rect 800 40600 39823 40728
rect 800 40464 39120 40600
rect 880 40320 39120 40464
rect 880 40184 39823 40320
rect 800 40056 39823 40184
rect 800 39776 39120 40056
rect 800 39648 39823 39776
rect 880 39368 39120 39648
rect 800 39240 39823 39368
rect 800 38960 39120 39240
rect 800 38832 39823 38960
rect 880 38552 39120 38832
rect 800 38288 39823 38552
rect 800 38016 39120 38288
rect 880 38008 39120 38016
rect 880 37880 39823 38008
rect 880 37736 39120 37880
rect 800 37600 39120 37736
rect 800 37472 39823 37600
rect 800 37200 39120 37472
rect 880 37192 39120 37200
rect 880 36928 39823 37192
rect 880 36920 39120 36928
rect 800 36648 39120 36920
rect 800 36520 39823 36648
rect 800 36384 39120 36520
rect 880 36240 39120 36384
rect 880 36112 39823 36240
rect 880 36104 39120 36112
rect 800 35832 39120 36104
rect 800 35568 39823 35832
rect 880 35288 39120 35568
rect 800 35160 39823 35288
rect 800 34880 39120 35160
rect 800 34752 39823 34880
rect 880 34472 39120 34752
rect 800 34344 39823 34472
rect 800 34064 39120 34344
rect 800 33936 39823 34064
rect 880 33800 39823 33936
rect 880 33656 39120 33800
rect 800 33520 39120 33656
rect 800 33392 39823 33520
rect 800 33256 39120 33392
rect 880 33112 39120 33256
rect 880 32984 39823 33112
rect 880 32976 39120 32984
rect 800 32704 39120 32976
rect 800 32440 39823 32704
rect 880 32160 39120 32440
rect 800 32032 39823 32160
rect 800 31752 39120 32032
rect 800 31624 39823 31752
rect 880 31344 39120 31624
rect 800 31216 39823 31344
rect 800 30936 39120 31216
rect 800 30808 39823 30936
rect 880 30672 39823 30808
rect 880 30528 39120 30672
rect 800 30392 39120 30528
rect 800 30264 39823 30392
rect 800 29992 39120 30264
rect 880 29984 39120 29992
rect 880 29856 39823 29984
rect 880 29712 39120 29856
rect 800 29576 39120 29712
rect 800 29312 39823 29576
rect 800 29176 39120 29312
rect 880 29032 39120 29176
rect 880 28904 39823 29032
rect 880 28896 39120 28904
rect 800 28624 39120 28896
rect 800 28496 39823 28624
rect 800 28360 39120 28496
rect 880 28216 39120 28360
rect 880 28088 39823 28216
rect 880 28080 39120 28088
rect 800 27808 39120 28080
rect 800 27544 39823 27808
rect 880 27264 39120 27544
rect 800 27136 39823 27264
rect 800 26864 39120 27136
rect 880 26856 39120 26864
rect 880 26728 39823 26856
rect 880 26584 39120 26728
rect 800 26448 39120 26584
rect 800 26184 39823 26448
rect 800 26048 39120 26184
rect 880 25904 39120 26048
rect 880 25776 39823 25904
rect 880 25768 39120 25776
rect 800 25496 39120 25768
rect 800 25368 39823 25496
rect 800 25232 39120 25368
rect 880 25088 39120 25232
rect 880 24960 39823 25088
rect 880 24952 39120 24960
rect 800 24680 39120 24952
rect 800 24416 39823 24680
rect 880 24136 39120 24416
rect 800 24008 39823 24136
rect 800 23728 39120 24008
rect 800 23600 39823 23728
rect 880 23320 39120 23600
rect 800 23056 39823 23320
rect 800 22784 39120 23056
rect 880 22776 39120 22784
rect 880 22648 39823 22776
rect 880 22504 39120 22648
rect 800 22368 39120 22504
rect 800 22240 39823 22368
rect 800 21968 39120 22240
rect 880 21960 39120 21968
rect 880 21696 39823 21960
rect 880 21688 39120 21696
rect 800 21416 39120 21688
rect 800 21288 39823 21416
rect 800 21152 39120 21288
rect 880 21008 39120 21152
rect 880 20880 39823 21008
rect 880 20872 39120 20880
rect 800 20600 39120 20872
rect 800 20472 39823 20600
rect 880 20192 39120 20472
rect 800 19928 39823 20192
rect 800 19656 39120 19928
rect 880 19648 39120 19656
rect 880 19520 39823 19648
rect 880 19376 39120 19520
rect 800 19240 39120 19376
rect 800 19112 39823 19240
rect 800 18840 39120 19112
rect 880 18832 39120 18840
rect 880 18568 39823 18832
rect 880 18560 39120 18568
rect 800 18288 39120 18560
rect 800 18160 39823 18288
rect 800 18024 39120 18160
rect 880 17880 39120 18024
rect 880 17752 39823 17880
rect 880 17744 39120 17752
rect 800 17472 39120 17744
rect 800 17344 39823 17472
rect 800 17208 39120 17344
rect 880 17064 39120 17208
rect 880 16928 39823 17064
rect 800 16800 39823 16928
rect 800 16520 39120 16800
rect 800 16392 39823 16520
rect 880 16112 39120 16392
rect 800 15984 39823 16112
rect 800 15704 39120 15984
rect 800 15576 39823 15704
rect 880 15440 39823 15576
rect 880 15296 39120 15440
rect 800 15160 39120 15296
rect 800 15032 39823 15160
rect 800 14760 39120 15032
rect 880 14752 39120 14760
rect 880 14624 39823 14752
rect 880 14480 39120 14624
rect 800 14344 39120 14480
rect 800 14216 39823 14344
rect 800 13944 39120 14216
rect 880 13936 39120 13944
rect 880 13672 39823 13936
rect 880 13664 39120 13672
rect 800 13392 39120 13664
rect 800 13264 39823 13392
rect 880 12984 39120 13264
rect 800 12856 39823 12984
rect 800 12576 39120 12856
rect 800 12448 39823 12576
rect 880 12312 39823 12448
rect 880 12168 39120 12312
rect 800 12032 39120 12168
rect 800 11904 39823 12032
rect 800 11632 39120 11904
rect 880 11624 39120 11632
rect 880 11496 39823 11624
rect 880 11352 39120 11496
rect 800 11216 39120 11352
rect 800 10952 39823 11216
rect 800 10816 39120 10952
rect 880 10672 39120 10816
rect 880 10544 39823 10672
rect 880 10536 39120 10544
rect 800 10264 39120 10536
rect 800 10136 39823 10264
rect 800 10000 39120 10136
rect 880 9856 39120 10000
rect 880 9728 39823 9856
rect 880 9720 39120 9728
rect 800 9448 39120 9720
rect 800 9184 39823 9448
rect 880 8904 39120 9184
rect 800 8776 39823 8904
rect 800 8496 39120 8776
rect 800 8368 39823 8496
rect 880 8088 39120 8368
rect 800 7824 39823 8088
rect 800 7552 39120 7824
rect 880 7544 39120 7552
rect 880 7416 39823 7544
rect 880 7272 39120 7416
rect 800 7136 39120 7272
rect 800 7008 39823 7136
rect 800 6872 39120 7008
rect 880 6728 39120 6872
rect 880 6600 39823 6728
rect 880 6592 39120 6600
rect 800 6320 39120 6592
rect 800 6056 39823 6320
rect 880 5776 39120 6056
rect 800 5648 39823 5776
rect 800 5368 39120 5648
rect 800 5240 39823 5368
rect 880 4960 39120 5240
rect 800 4696 39823 4960
rect 800 4424 39120 4696
rect 880 4416 39120 4424
rect 880 4288 39823 4416
rect 880 4144 39120 4288
rect 800 4008 39120 4144
rect 800 3880 39823 4008
rect 800 3608 39120 3880
rect 880 3600 39120 3608
rect 880 3472 39823 3600
rect 880 3328 39120 3472
rect 800 3192 39120 3328
rect 800 2928 39823 3192
rect 800 2792 39120 2928
rect 880 2648 39120 2792
rect 880 2520 39823 2648
rect 880 2512 39120 2520
rect 800 2240 39120 2512
rect 800 2112 39823 2240
rect 800 1976 39120 2112
rect 880 1832 39120 1976
rect 880 1696 39823 1832
rect 800 1568 39823 1696
rect 800 1288 39120 1568
rect 800 1160 39823 1288
rect 880 880 39120 1160
rect 800 752 39823 880
rect 800 480 39120 752
rect 880 472 39120 480
rect 880 344 39823 472
rect 880 200 39120 344
rect 800 171 39120 200
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
<< labels >>
rlabel metal2 s 110 119200 166 120800 6 dsi[0]
port 1 nsew signal output
rlabel metal2 s 294 119200 350 120800 6 dsi[1]
port 2 nsew signal output
rlabel metal2 s 570 119200 626 120800 6 dsi[2]
port 3 nsew signal output
rlabel metal2 s 754 119200 810 120800 6 dsi[3]
port 4 nsew signal output
rlabel metal2 s 1030 119200 1086 120800 6 dsi[4]
port 5 nsew signal output
rlabel metal2 s 1214 119200 1270 120800 6 dsi[5]
port 6 nsew signal output
rlabel metal2 s 1490 119200 1546 120800 6 dsi[6]
port 7 nsew signal output
rlabel metal2 s 1674 119200 1730 120800 6 dsi[7]
port 8 nsew signal output
rlabel metal2 s 1950 119200 2006 120800 6 io_in[0]
port 9 nsew signal input
rlabel metal2 s 8850 119200 8906 120800 6 io_in[10]
port 10 nsew signal input
rlabel metal2 s 9586 119200 9642 120800 6 io_in[11]
port 11 nsew signal input
rlabel metal2 s 10230 119200 10286 120800 6 io_in[12]
port 12 nsew signal input
rlabel metal2 s 10966 119200 11022 120800 6 io_in[13]
port 13 nsew signal input
rlabel metal2 s 11610 119200 11666 120800 6 io_in[14]
port 14 nsew signal input
rlabel metal2 s 12346 119200 12402 120800 6 io_in[15]
port 15 nsew signal input
rlabel metal2 s 12990 119200 13046 120800 6 io_in[16]
port 16 nsew signal input
rlabel metal2 s 13726 119200 13782 120800 6 io_in[17]
port 17 nsew signal input
rlabel metal2 s 14370 119200 14426 120800 6 io_in[18]
port 18 nsew signal input
rlabel metal2 s 15106 119200 15162 120800 6 io_in[19]
port 19 nsew signal input
rlabel metal2 s 2594 119200 2650 120800 6 io_in[1]
port 20 nsew signal input
rlabel metal2 s 15750 119200 15806 120800 6 io_in[20]
port 21 nsew signal input
rlabel metal2 s 16486 119200 16542 120800 6 io_in[21]
port 22 nsew signal input
rlabel metal2 s 17222 119200 17278 120800 6 io_in[22]
port 23 nsew signal input
rlabel metal2 s 17866 119200 17922 120800 6 io_in[23]
port 24 nsew signal input
rlabel metal2 s 18602 119200 18658 120800 6 io_in[24]
port 25 nsew signal input
rlabel metal2 s 19246 119200 19302 120800 6 io_in[25]
port 26 nsew signal input
rlabel metal2 s 19982 119200 20038 120800 6 io_in[26]
port 27 nsew signal input
rlabel metal2 s 20626 119200 20682 120800 6 io_in[27]
port 28 nsew signal input
rlabel metal2 s 21362 119200 21418 120800 6 io_in[28]
port 29 nsew signal input
rlabel metal2 s 22006 119200 22062 120800 6 io_in[29]
port 30 nsew signal input
rlabel metal2 s 3330 119200 3386 120800 6 io_in[2]
port 31 nsew signal input
rlabel metal2 s 22742 119200 22798 120800 6 io_in[30]
port 32 nsew signal input
rlabel metal2 s 23386 119200 23442 120800 6 io_in[31]
port 33 nsew signal input
rlabel metal2 s 24122 119200 24178 120800 6 io_in[32]
port 34 nsew signal input
rlabel metal2 s 24858 119200 24914 120800 6 io_in[33]
port 35 nsew signal input
rlabel metal2 s 25502 119200 25558 120800 6 io_in[34]
port 36 nsew signal input
rlabel metal2 s 26238 119200 26294 120800 6 io_in[35]
port 37 nsew signal input
rlabel metal2 s 26882 119200 26938 120800 6 io_in[36]
port 38 nsew signal input
rlabel metal2 s 27618 119200 27674 120800 6 io_in[37]
port 39 nsew signal input
rlabel metal2 s 3974 119200 4030 120800 6 io_in[3]
port 40 nsew signal input
rlabel metal2 s 4710 119200 4766 120800 6 io_in[4]
port 41 nsew signal input
rlabel metal2 s 5354 119200 5410 120800 6 io_in[5]
port 42 nsew signal input
rlabel metal2 s 6090 119200 6146 120800 6 io_in[6]
port 43 nsew signal input
rlabel metal2 s 6734 119200 6790 120800 6 io_in[7]
port 44 nsew signal input
rlabel metal2 s 7470 119200 7526 120800 6 io_in[8]
port 45 nsew signal input
rlabel metal2 s 8206 119200 8262 120800 6 io_in[9]
port 46 nsew signal input
rlabel metal2 s 2134 119200 2190 120800 6 io_oeb[0]
port 47 nsew signal output
rlabel metal2 s 9126 119200 9182 120800 6 io_oeb[10]
port 48 nsew signal output
rlabel metal2 s 9770 119200 9826 120800 6 io_oeb[11]
port 49 nsew signal output
rlabel metal2 s 10506 119200 10562 120800 6 io_oeb[12]
port 50 nsew signal output
rlabel metal2 s 11150 119200 11206 120800 6 io_oeb[13]
port 51 nsew signal output
rlabel metal2 s 11886 119200 11942 120800 6 io_oeb[14]
port 52 nsew signal output
rlabel metal2 s 12530 119200 12586 120800 6 io_oeb[15]
port 53 nsew signal output
rlabel metal2 s 13266 119200 13322 120800 6 io_oeb[16]
port 54 nsew signal output
rlabel metal2 s 13910 119200 13966 120800 6 io_oeb[17]
port 55 nsew signal output
rlabel metal2 s 14646 119200 14702 120800 6 io_oeb[18]
port 56 nsew signal output
rlabel metal2 s 15290 119200 15346 120800 6 io_oeb[19]
port 57 nsew signal output
rlabel metal2 s 2870 119200 2926 120800 6 io_oeb[1]
port 58 nsew signal output
rlabel metal2 s 16026 119200 16082 120800 6 io_oeb[20]
port 59 nsew signal output
rlabel metal2 s 16762 119200 16818 120800 6 io_oeb[21]
port 60 nsew signal output
rlabel metal2 s 17406 119200 17462 120800 6 io_oeb[22]
port 61 nsew signal output
rlabel metal2 s 18142 119200 18198 120800 6 io_oeb[23]
port 62 nsew signal output
rlabel metal2 s 18786 119200 18842 120800 6 io_oeb[24]
port 63 nsew signal output
rlabel metal2 s 19522 119200 19578 120800 6 io_oeb[25]
port 64 nsew signal output
rlabel metal2 s 20166 119200 20222 120800 6 io_oeb[26]
port 65 nsew signal output
rlabel metal2 s 20902 119200 20958 120800 6 io_oeb[27]
port 66 nsew signal output
rlabel metal2 s 21546 119200 21602 120800 6 io_oeb[28]
port 67 nsew signal output
rlabel metal2 s 22282 119200 22338 120800 6 io_oeb[29]
port 68 nsew signal output
rlabel metal2 s 3514 119200 3570 120800 6 io_oeb[2]
port 69 nsew signal output
rlabel metal2 s 22926 119200 22982 120800 6 io_oeb[30]
port 70 nsew signal output
rlabel metal2 s 23662 119200 23718 120800 6 io_oeb[31]
port 71 nsew signal output
rlabel metal2 s 24398 119200 24454 120800 6 io_oeb[32]
port 72 nsew signal output
rlabel metal2 s 25042 119200 25098 120800 6 io_oeb[33]
port 73 nsew signal output
rlabel metal2 s 25778 119200 25834 120800 6 io_oeb[34]
port 74 nsew signal output
rlabel metal2 s 26422 119200 26478 120800 6 io_oeb[35]
port 75 nsew signal output
rlabel metal2 s 27158 119200 27214 120800 6 io_oeb[36]
port 76 nsew signal output
rlabel metal2 s 27802 119200 27858 120800 6 io_oeb[37]
port 77 nsew signal output
rlabel metal2 s 4250 119200 4306 120800 6 io_oeb[3]
port 78 nsew signal output
rlabel metal2 s 4894 119200 4950 120800 6 io_oeb[4]
port 79 nsew signal output
rlabel metal2 s 5630 119200 5686 120800 6 io_oeb[5]
port 80 nsew signal output
rlabel metal2 s 6274 119200 6330 120800 6 io_oeb[6]
port 81 nsew signal output
rlabel metal2 s 7010 119200 7066 120800 6 io_oeb[7]
port 82 nsew signal output
rlabel metal2 s 7654 119200 7710 120800 6 io_oeb[8]
port 83 nsew signal output
rlabel metal2 s 8390 119200 8446 120800 6 io_oeb[9]
port 84 nsew signal output
rlabel metal2 s 2410 119200 2466 120800 6 io_out[0]
port 85 nsew signal output
rlabel metal2 s 9310 119200 9366 120800 6 io_out[10]
port 86 nsew signal output
rlabel metal2 s 10046 119200 10102 120800 6 io_out[11]
port 87 nsew signal output
rlabel metal2 s 10690 119200 10746 120800 6 io_out[12]
port 88 nsew signal output
rlabel metal2 s 11426 119200 11482 120800 6 io_out[13]
port 89 nsew signal output
rlabel metal2 s 12070 119200 12126 120800 6 io_out[14]
port 90 nsew signal output
rlabel metal2 s 12806 119200 12862 120800 6 io_out[15]
port 91 nsew signal output
rlabel metal2 s 13450 119200 13506 120800 6 io_out[16]
port 92 nsew signal output
rlabel metal2 s 14186 119200 14242 120800 6 io_out[17]
port 93 nsew signal output
rlabel metal2 s 14830 119200 14886 120800 6 io_out[18]
port 94 nsew signal output
rlabel metal2 s 15566 119200 15622 120800 6 io_out[19]
port 95 nsew signal output
rlabel metal2 s 3054 119200 3110 120800 6 io_out[1]
port 96 nsew signal output
rlabel metal2 s 16302 119200 16358 120800 6 io_out[20]
port 97 nsew signal output
rlabel metal2 s 16946 119200 17002 120800 6 io_out[21]
port 98 nsew signal output
rlabel metal2 s 17682 119200 17738 120800 6 io_out[22]
port 99 nsew signal output
rlabel metal2 s 18326 119200 18382 120800 6 io_out[23]
port 100 nsew signal output
rlabel metal2 s 19062 119200 19118 120800 6 io_out[24]
port 101 nsew signal output
rlabel metal2 s 19706 119200 19762 120800 6 io_out[25]
port 102 nsew signal output
rlabel metal2 s 20442 119200 20498 120800 6 io_out[26]
port 103 nsew signal output
rlabel metal2 s 21086 119200 21142 120800 6 io_out[27]
port 104 nsew signal output
rlabel metal2 s 21822 119200 21878 120800 6 io_out[28]
port 105 nsew signal output
rlabel metal2 s 22466 119200 22522 120800 6 io_out[29]
port 106 nsew signal output
rlabel metal2 s 3790 119200 3846 120800 6 io_out[2]
port 107 nsew signal output
rlabel metal2 s 23202 119200 23258 120800 6 io_out[30]
port 108 nsew signal output
rlabel metal2 s 23846 119200 23902 120800 6 io_out[31]
port 109 nsew signal output
rlabel metal2 s 24582 119200 24638 120800 6 io_out[32]
port 110 nsew signal output
rlabel metal2 s 25318 119200 25374 120800 6 io_out[33]
port 111 nsew signal output
rlabel metal2 s 25962 119200 26018 120800 6 io_out[34]
port 112 nsew signal output
rlabel metal2 s 26698 119200 26754 120800 6 io_out[35]
port 113 nsew signal output
rlabel metal2 s 27342 119200 27398 120800 6 io_out[36]
port 114 nsew signal output
rlabel metal2 s 28078 119200 28134 120800 6 io_out[37]
port 115 nsew signal output
rlabel metal2 s 4434 119200 4490 120800 6 io_out[3]
port 116 nsew signal output
rlabel metal2 s 5170 119200 5226 120800 6 io_out[4]
port 117 nsew signal output
rlabel metal2 s 5814 119200 5870 120800 6 io_out[5]
port 118 nsew signal output
rlabel metal2 s 6550 119200 6606 120800 6 io_out[6]
port 119 nsew signal output
rlabel metal2 s 7194 119200 7250 120800 6 io_out[7]
port 120 nsew signal output
rlabel metal2 s 7930 119200 7986 120800 6 io_out[8]
port 121 nsew signal output
rlabel metal2 s 8666 119200 8722 120800 6 io_out[9]
port 122 nsew signal output
rlabel metal2 s 754 -800 810 800 8 irq[0]
port 123 nsew signal output
rlabel metal2 s 1030 -800 1086 800 8 irq[1]
port 124 nsew signal output
rlabel metal2 s 1398 -800 1454 800 8 irq[2]
port 125 nsew signal output
rlabel metal2 s 31942 119200 31998 120800 6 m_irqs[0]
port 126 nsew signal input
rlabel metal2 s 34334 119200 34390 120800 6 m_irqs[10]
port 127 nsew signal input
rlabel metal2 s 34518 119200 34574 120800 6 m_irqs[11]
port 128 nsew signal input
rlabel metal2 s 32218 119200 32274 120800 6 m_irqs[1]
port 129 nsew signal input
rlabel metal2 s 32494 119200 32550 120800 6 m_irqs[2]
port 130 nsew signal input
rlabel metal2 s 32678 119200 32734 120800 6 m_irqs[3]
port 131 nsew signal input
rlabel metal2 s 32954 119200 33010 120800 6 m_irqs[4]
port 132 nsew signal input
rlabel metal2 s 33138 119200 33194 120800 6 m_irqs[5]
port 133 nsew signal input
rlabel metal2 s 33414 119200 33470 120800 6 m_irqs[6]
port 134 nsew signal input
rlabel metal2 s 33598 119200 33654 120800 6 m_irqs[7]
port 135 nsew signal input
rlabel metal2 s 33874 119200 33930 120800 6 m_irqs[8]
port 136 nsew signal input
rlabel metal2 s 34058 119200 34114 120800 6 m_irqs[9]
port 137 nsew signal input
rlabel metal2 s 35530 -800 35586 800 8 m_wb_clk_i
port 138 nsew signal output
rlabel metal2 s 34794 119200 34850 120800 6 m_wb_rst_i
port 139 nsew signal output
rlabel metal2 s 35898 -800 35954 800 8 m_wbs_ack_o[0]
port 140 nsew signal input
rlabel metal3 s -800 113704 800 113824 4 m_wbs_ack_o[10]
port 141 nsew signal input
rlabel metal2 s 38474 119200 38530 120800 6 m_wbs_ack_o[11]
port 142 nsew signal input
rlabel metal3 s -800 104184 800 104304 4 m_wbs_ack_o[1]
port 143 nsew signal input
rlabel metal3 s -800 105816 800 105936 4 m_wbs_ack_o[2]
port 144 nsew signal input
rlabel metal2 s 35438 119200 35494 120800 6 m_wbs_ack_o[3]
port 145 nsew signal input
rlabel metal3 s -800 108944 800 109064 4 m_wbs_ack_o[4]
port 146 nsew signal input
rlabel metal2 s 36358 119200 36414 120800 6 m_wbs_ack_o[5]
port 147 nsew signal input
rlabel metal2 s 37094 119200 37150 120800 6 m_wbs_ack_o[6]
port 148 nsew signal input
rlabel metal2 s 37554 119200 37610 120800 6 m_wbs_ack_o[7]
port 149 nsew signal input
rlabel metal3 s 39200 116016 40800 116136 6 m_wbs_ack_o[8]
port 150 nsew signal input
rlabel metal2 s 37462 -800 37518 800 8 m_wbs_ack_o[9]
port 151 nsew signal input
rlabel metal3 s -800 103368 800 103488 4 m_wbs_adr_i[0]
port 152 nsew signal output
rlabel metal3 s -800 114520 800 114640 4 m_wbs_adr_i[10]
port 153 nsew signal output
rlabel metal2 s 38106 -800 38162 800 8 m_wbs_adr_i[11]
port 154 nsew signal output
rlabel metal2 s 36542 -800 36598 800 8 m_wbs_adr_i[1]
port 155 nsew signal output
rlabel metal3 s -800 106632 800 106752 4 m_wbs_adr_i[2]
port 156 nsew signal output
rlabel metal3 s -800 108128 800 108248 4 m_wbs_adr_i[3]
port 157 nsew signal output
rlabel metal3 s -800 109760 800 109880 4 m_wbs_adr_i[4]
port 158 nsew signal output
rlabel metal2 s 36634 119200 36690 120800 6 m_wbs_adr_i[5]
port 159 nsew signal output
rlabel metal3 s -800 110576 800 110696 4 m_wbs_adr_i[6]
port 160 nsew signal output
rlabel metal3 s 39200 115064 40800 115184 6 m_wbs_adr_i[7]
port 161 nsew signal output
rlabel metal2 s 38014 119200 38070 120800 6 m_wbs_adr_i[8]
port 162 nsew signal output
rlabel metal3 s -800 113024 800 113144 4 m_wbs_adr_i[9]
port 163 nsew signal output
rlabel metal2 s 36174 -800 36230 800 8 m_wbs_cs_i[0]
port 164 nsew signal output
rlabel metal2 s 38198 119200 38254 120800 6 m_wbs_cs_i[10]
port 165 nsew signal output
rlabel metal2 s 38474 -800 38530 800 8 m_wbs_cs_i[11]
port 166 nsew signal output
rlabel metal2 s 35254 119200 35310 120800 6 m_wbs_cs_i[1]
port 167 nsew signal output
rlabel metal3 s 39200 114656 40800 114776 6 m_wbs_cs_i[2]
port 168 nsew signal output
rlabel metal2 s 35714 119200 35770 120800 6 m_wbs_cs_i[3]
port 169 nsew signal output
rlabel metal2 s 36174 119200 36230 120800 6 m_wbs_cs_i[4]
port 170 nsew signal output
rlabel metal2 s 36818 119200 36874 120800 6 m_wbs_cs_i[5]
port 171 nsew signal output
rlabel metal2 s 37278 119200 37334 120800 6 m_wbs_cs_i[6]
port 172 nsew signal output
rlabel metal2 s 37738 119200 37794 120800 6 m_wbs_cs_i[7]
port 173 nsew signal output
rlabel metal3 s 39200 116424 40800 116544 6 m_wbs_cs_i[8]
port 174 nsew signal output
rlabel metal3 s 39200 116832 40800 116952 6 m_wbs_cs_i[9]
port 175 nsew signal output
rlabel metal2 s 34978 119200 35034 120800 6 m_wbs_dat_i[0]
port 176 nsew signal output
rlabel metal2 s 37830 -800 37886 800 8 m_wbs_dat_i[10]
port 177 nsew signal output
rlabel metal3 s -800 115336 800 115456 4 m_wbs_dat_i[11]
port 178 nsew signal output
rlabel metal2 s 38658 119200 38714 120800 6 m_wbs_dat_i[12]
port 179 nsew signal output
rlabel metal3 s 39200 117784 40800 117904 6 m_wbs_dat_i[13]
port 180 nsew signal output
rlabel metal3 s -800 116152 800 116272 4 m_wbs_dat_i[14]
port 181 nsew signal output
rlabel metal2 s 38934 119200 38990 120800 6 m_wbs_dat_i[15]
port 182 nsew signal output
rlabel metal3 s -800 116968 800 117088 4 m_wbs_dat_i[16]
port 183 nsew signal output
rlabel metal3 s 39200 118192 40800 118312 6 m_wbs_dat_i[17]
port 184 nsew signal output
rlabel metal3 s 39200 118736 40800 118856 6 m_wbs_dat_i[18]
port 185 nsew signal output
rlabel metal2 s 38750 -800 38806 800 8 m_wbs_dat_i[19]
port 186 nsew signal output
rlabel metal3 s -800 105000 800 105120 4 m_wbs_dat_i[1]
port 187 nsew signal output
rlabel metal2 s 39118 -800 39174 800 8 m_wbs_dat_i[20]
port 188 nsew signal output
rlabel metal2 s 39118 119200 39174 120800 6 m_wbs_dat_i[21]
port 189 nsew signal output
rlabel metal3 s -800 117784 800 117904 4 m_wbs_dat_i[22]
port 190 nsew signal output
rlabel metal2 s 39394 119200 39450 120800 6 m_wbs_dat_i[23]
port 191 nsew signal output
rlabel metal2 s 39578 119200 39634 120800 6 m_wbs_dat_i[24]
port 192 nsew signal output
rlabel metal2 s 39394 -800 39450 800 8 m_wbs_dat_i[25]
port 193 nsew signal output
rlabel metal3 s -800 118600 800 118720 4 m_wbs_dat_i[26]
port 194 nsew signal output
rlabel metal3 s -800 119416 800 119536 4 m_wbs_dat_i[27]
port 195 nsew signal output
rlabel metal2 s 39762 -800 39818 800 8 m_wbs_dat_i[28]
port 196 nsew signal output
rlabel metal3 s 39200 119144 40800 119264 6 m_wbs_dat_i[29]
port 197 nsew signal output
rlabel metal3 s -800 107312 800 107432 4 m_wbs_dat_i[2]
port 198 nsew signal output
rlabel metal3 s 39200 119552 40800 119672 6 m_wbs_dat_i[30]
port 199 nsew signal output
rlabel metal2 s 39854 119200 39910 120800 6 m_wbs_dat_i[31]
port 200 nsew signal output
rlabel metal2 s 35898 119200 35954 120800 6 m_wbs_dat_i[3]
port 201 nsew signal output
rlabel metal2 s 36818 -800 36874 800 8 m_wbs_dat_i[4]
port 202 nsew signal output
rlabel metal2 s 37186 -800 37242 800 8 m_wbs_dat_i[5]
port 203 nsew signal output
rlabel metal3 s -800 111392 800 111512 4 m_wbs_dat_i[6]
port 204 nsew signal output
rlabel metal3 s 39200 115608 40800 115728 6 m_wbs_dat_i[7]
port 205 nsew signal output
rlabel metal3 s -800 112208 800 112328 4 m_wbs_dat_i[8]
port 206 nsew signal output
rlabel metal3 s 39200 117376 40800 117496 6 m_wbs_dat_i[9]
port 207 nsew signal output
rlabel metal3 s 39200 144 40800 264 6 m_wbs_dat_o_0[0]
port 208 nsew signal input
rlabel metal3 s 39200 4496 40800 4616 6 m_wbs_dat_o_0[10]
port 209 nsew signal input
rlabel metal3 s 39200 5040 40800 5160 6 m_wbs_dat_o_0[11]
port 210 nsew signal input
rlabel metal3 s 39200 5448 40800 5568 6 m_wbs_dat_o_0[12]
port 211 nsew signal input
rlabel metal3 s 39200 5856 40800 5976 6 m_wbs_dat_o_0[13]
port 212 nsew signal input
rlabel metal3 s 39200 6400 40800 6520 6 m_wbs_dat_o_0[14]
port 213 nsew signal input
rlabel metal3 s 39200 6808 40800 6928 6 m_wbs_dat_o_0[15]
port 214 nsew signal input
rlabel metal3 s 39200 7216 40800 7336 6 m_wbs_dat_o_0[16]
port 215 nsew signal input
rlabel metal3 s 39200 7624 40800 7744 6 m_wbs_dat_o_0[17]
port 216 nsew signal input
rlabel metal3 s 39200 8168 40800 8288 6 m_wbs_dat_o_0[18]
port 217 nsew signal input
rlabel metal3 s 39200 8576 40800 8696 6 m_wbs_dat_o_0[19]
port 218 nsew signal input
rlabel metal3 s 39200 552 40800 672 6 m_wbs_dat_o_0[1]
port 219 nsew signal input
rlabel metal3 s 39200 8984 40800 9104 6 m_wbs_dat_o_0[20]
port 220 nsew signal input
rlabel metal3 s 39200 9528 40800 9648 6 m_wbs_dat_o_0[21]
port 221 nsew signal input
rlabel metal3 s 39200 9936 40800 10056 6 m_wbs_dat_o_0[22]
port 222 nsew signal input
rlabel metal3 s 39200 10344 40800 10464 6 m_wbs_dat_o_0[23]
port 223 nsew signal input
rlabel metal3 s 39200 10752 40800 10872 6 m_wbs_dat_o_0[24]
port 224 nsew signal input
rlabel metal3 s 39200 11296 40800 11416 6 m_wbs_dat_o_0[25]
port 225 nsew signal input
rlabel metal3 s 39200 11704 40800 11824 6 m_wbs_dat_o_0[26]
port 226 nsew signal input
rlabel metal3 s 39200 12112 40800 12232 6 m_wbs_dat_o_0[27]
port 227 nsew signal input
rlabel metal3 s 39200 12656 40800 12776 6 m_wbs_dat_o_0[28]
port 228 nsew signal input
rlabel metal3 s 39200 13064 40800 13184 6 m_wbs_dat_o_0[29]
port 229 nsew signal input
rlabel metal3 s 39200 960 40800 1080 6 m_wbs_dat_o_0[2]
port 230 nsew signal input
rlabel metal3 s 39200 13472 40800 13592 6 m_wbs_dat_o_0[30]
port 231 nsew signal input
rlabel metal3 s 39200 14016 40800 14136 6 m_wbs_dat_o_0[31]
port 232 nsew signal input
rlabel metal3 s 39200 1368 40800 1488 6 m_wbs_dat_o_0[3]
port 233 nsew signal input
rlabel metal3 s 39200 1912 40800 2032 6 m_wbs_dat_o_0[4]
port 234 nsew signal input
rlabel metal3 s 39200 2320 40800 2440 6 m_wbs_dat_o_0[5]
port 235 nsew signal input
rlabel metal3 s 39200 2728 40800 2848 6 m_wbs_dat_o_0[6]
port 236 nsew signal input
rlabel metal3 s 39200 3272 40800 3392 6 m_wbs_dat_o_0[7]
port 237 nsew signal input
rlabel metal3 s 39200 3680 40800 3800 6 m_wbs_dat_o_0[8]
port 238 nsew signal input
rlabel metal3 s 39200 4088 40800 4208 6 m_wbs_dat_o_0[9]
port 239 nsew signal input
rlabel metal3 s 39200 14832 40800 14952 6 m_wbs_dat_o_10[0]
port 240 nsew signal input
rlabel metal3 s 39200 28296 40800 28416 6 m_wbs_dat_o_10[10]
port 241 nsew signal input
rlabel metal3 s 39200 29656 40800 29776 6 m_wbs_dat_o_10[11]
port 242 nsew signal input
rlabel metal3 s 39200 31016 40800 31136 6 m_wbs_dat_o_10[12]
port 243 nsew signal input
rlabel metal3 s 39200 32240 40800 32360 6 m_wbs_dat_o_10[13]
port 244 nsew signal input
rlabel metal3 s 39200 33600 40800 33720 6 m_wbs_dat_o_10[14]
port 245 nsew signal input
rlabel metal3 s 39200 34960 40800 35080 6 m_wbs_dat_o_10[15]
port 246 nsew signal input
rlabel metal3 s 39200 36320 40800 36440 6 m_wbs_dat_o_10[16]
port 247 nsew signal input
rlabel metal3 s 39200 37680 40800 37800 6 m_wbs_dat_o_10[17]
port 248 nsew signal input
rlabel metal3 s 39200 39040 40800 39160 6 m_wbs_dat_o_10[18]
port 249 nsew signal input
rlabel metal3 s 39200 40400 40800 40520 6 m_wbs_dat_o_10[19]
port 250 nsew signal input
rlabel metal3 s 39200 16192 40800 16312 6 m_wbs_dat_o_10[1]
port 251 nsew signal input
rlabel metal3 s 39200 41760 40800 41880 6 m_wbs_dat_o_10[20]
port 252 nsew signal input
rlabel metal3 s 39200 42984 40800 43104 6 m_wbs_dat_o_10[21]
port 253 nsew signal input
rlabel metal3 s 39200 44344 40800 44464 6 m_wbs_dat_o_10[22]
port 254 nsew signal input
rlabel metal3 s 39200 45704 40800 45824 6 m_wbs_dat_o_10[23]
port 255 nsew signal input
rlabel metal3 s 39200 47064 40800 47184 6 m_wbs_dat_o_10[24]
port 256 nsew signal input
rlabel metal3 s 39200 48424 40800 48544 6 m_wbs_dat_o_10[25]
port 257 nsew signal input
rlabel metal3 s 39200 49784 40800 49904 6 m_wbs_dat_o_10[26]
port 258 nsew signal input
rlabel metal3 s 39200 51144 40800 51264 6 m_wbs_dat_o_10[27]
port 259 nsew signal input
rlabel metal3 s 39200 52504 40800 52624 6 m_wbs_dat_o_10[28]
port 260 nsew signal input
rlabel metal3 s 39200 53728 40800 53848 6 m_wbs_dat_o_10[29]
port 261 nsew signal input
rlabel metal3 s 39200 17552 40800 17672 6 m_wbs_dat_o_10[2]
port 262 nsew signal input
rlabel metal3 s 39200 55088 40800 55208 6 m_wbs_dat_o_10[30]
port 263 nsew signal input
rlabel metal3 s 39200 56448 40800 56568 6 m_wbs_dat_o_10[31]
port 264 nsew signal input
rlabel metal3 s 39200 18912 40800 19032 6 m_wbs_dat_o_10[3]
port 265 nsew signal input
rlabel metal3 s 39200 20272 40800 20392 6 m_wbs_dat_o_10[4]
port 266 nsew signal input
rlabel metal3 s 39200 21496 40800 21616 6 m_wbs_dat_o_10[5]
port 267 nsew signal input
rlabel metal3 s 39200 22856 40800 22976 6 m_wbs_dat_o_10[6]
port 268 nsew signal input
rlabel metal3 s 39200 24216 40800 24336 6 m_wbs_dat_o_10[7]
port 269 nsew signal input
rlabel metal3 s 39200 25576 40800 25696 6 m_wbs_dat_o_10[8]
port 270 nsew signal input
rlabel metal3 s 39200 26936 40800 27056 6 m_wbs_dat_o_10[9]
port 271 nsew signal input
rlabel metal3 s 39200 15240 40800 15360 6 m_wbs_dat_o_11[0]
port 272 nsew signal input
rlabel metal3 s 39200 28704 40800 28824 6 m_wbs_dat_o_11[10]
port 273 nsew signal input
rlabel metal3 s 39200 30064 40800 30184 6 m_wbs_dat_o_11[11]
port 274 nsew signal input
rlabel metal3 s 39200 31424 40800 31544 6 m_wbs_dat_o_11[12]
port 275 nsew signal input
rlabel metal3 s 39200 32784 40800 32904 6 m_wbs_dat_o_11[13]
port 276 nsew signal input
rlabel metal3 s 39200 34144 40800 34264 6 m_wbs_dat_o_11[14]
port 277 nsew signal input
rlabel metal3 s 39200 35368 40800 35488 6 m_wbs_dat_o_11[15]
port 278 nsew signal input
rlabel metal3 s 39200 36728 40800 36848 6 m_wbs_dat_o_11[16]
port 279 nsew signal input
rlabel metal3 s 39200 38088 40800 38208 6 m_wbs_dat_o_11[17]
port 280 nsew signal input
rlabel metal3 s 39200 39448 40800 39568 6 m_wbs_dat_o_11[18]
port 281 nsew signal input
rlabel metal3 s 39200 40808 40800 40928 6 m_wbs_dat_o_11[19]
port 282 nsew signal input
rlabel metal3 s 39200 16600 40800 16720 6 m_wbs_dat_o_11[1]
port 283 nsew signal input
rlabel metal3 s 39200 42168 40800 42288 6 m_wbs_dat_o_11[20]
port 284 nsew signal input
rlabel metal3 s 39200 43528 40800 43648 6 m_wbs_dat_o_11[21]
port 285 nsew signal input
rlabel metal3 s 39200 44888 40800 45008 6 m_wbs_dat_o_11[22]
port 286 nsew signal input
rlabel metal3 s 39200 46112 40800 46232 6 m_wbs_dat_o_11[23]
port 287 nsew signal input
rlabel metal3 s 39200 47472 40800 47592 6 m_wbs_dat_o_11[24]
port 288 nsew signal input
rlabel metal3 s 39200 48832 40800 48952 6 m_wbs_dat_o_11[25]
port 289 nsew signal input
rlabel metal3 s 39200 50192 40800 50312 6 m_wbs_dat_o_11[26]
port 290 nsew signal input
rlabel metal3 s 39200 51552 40800 51672 6 m_wbs_dat_o_11[27]
port 291 nsew signal input
rlabel metal3 s 39200 52912 40800 53032 6 m_wbs_dat_o_11[28]
port 292 nsew signal input
rlabel metal3 s 39200 54272 40800 54392 6 m_wbs_dat_o_11[29]
port 293 nsew signal input
rlabel metal3 s 39200 17960 40800 18080 6 m_wbs_dat_o_11[2]
port 294 nsew signal input
rlabel metal3 s 39200 55632 40800 55752 6 m_wbs_dat_o_11[30]
port 295 nsew signal input
rlabel metal3 s 39200 56856 40800 56976 6 m_wbs_dat_o_11[31]
port 296 nsew signal input
rlabel metal3 s 39200 19320 40800 19440 6 m_wbs_dat_o_11[3]
port 297 nsew signal input
rlabel metal3 s 39200 20680 40800 20800 6 m_wbs_dat_o_11[4]
port 298 nsew signal input
rlabel metal3 s 39200 22040 40800 22160 6 m_wbs_dat_o_11[5]
port 299 nsew signal input
rlabel metal3 s 39200 23400 40800 23520 6 m_wbs_dat_o_11[6]
port 300 nsew signal input
rlabel metal3 s 39200 24760 40800 24880 6 m_wbs_dat_o_11[7]
port 301 nsew signal input
rlabel metal3 s 39200 25984 40800 26104 6 m_wbs_dat_o_11[8]
port 302 nsew signal input
rlabel metal3 s 39200 27344 40800 27464 6 m_wbs_dat_o_11[9]
port 303 nsew signal input
rlabel metal3 s 39200 14424 40800 14544 6 m_wbs_dat_o_1[0]
port 304 nsew signal input
rlabel metal3 s 39200 27888 40800 28008 6 m_wbs_dat_o_1[10]
port 305 nsew signal input
rlabel metal3 s 39200 29112 40800 29232 6 m_wbs_dat_o_1[11]
port 306 nsew signal input
rlabel metal3 s 39200 30472 40800 30592 6 m_wbs_dat_o_1[12]
port 307 nsew signal input
rlabel metal3 s 39200 31832 40800 31952 6 m_wbs_dat_o_1[13]
port 308 nsew signal input
rlabel metal3 s 39200 33192 40800 33312 6 m_wbs_dat_o_1[14]
port 309 nsew signal input
rlabel metal3 s 39200 34552 40800 34672 6 m_wbs_dat_o_1[15]
port 310 nsew signal input
rlabel metal3 s 39200 35912 40800 36032 6 m_wbs_dat_o_1[16]
port 311 nsew signal input
rlabel metal3 s 39200 37272 40800 37392 6 m_wbs_dat_o_1[17]
port 312 nsew signal input
rlabel metal3 s 39200 38632 40800 38752 6 m_wbs_dat_o_1[18]
port 313 nsew signal input
rlabel metal3 s 39200 39856 40800 39976 6 m_wbs_dat_o_1[19]
port 314 nsew signal input
rlabel metal3 s 39200 15784 40800 15904 6 m_wbs_dat_o_1[1]
port 315 nsew signal input
rlabel metal3 s 39200 41216 40800 41336 6 m_wbs_dat_o_1[20]
port 316 nsew signal input
rlabel metal3 s 39200 42576 40800 42696 6 m_wbs_dat_o_1[21]
port 317 nsew signal input
rlabel metal3 s 39200 43936 40800 44056 6 m_wbs_dat_o_1[22]
port 318 nsew signal input
rlabel metal3 s 39200 45296 40800 45416 6 m_wbs_dat_o_1[23]
port 319 nsew signal input
rlabel metal3 s 39200 46656 40800 46776 6 m_wbs_dat_o_1[24]
port 320 nsew signal input
rlabel metal3 s 39200 48016 40800 48136 6 m_wbs_dat_o_1[25]
port 321 nsew signal input
rlabel metal3 s 39200 49376 40800 49496 6 m_wbs_dat_o_1[26]
port 322 nsew signal input
rlabel metal3 s 39200 50600 40800 50720 6 m_wbs_dat_o_1[27]
port 323 nsew signal input
rlabel metal3 s 39200 51960 40800 52080 6 m_wbs_dat_o_1[28]
port 324 nsew signal input
rlabel metal3 s 39200 53320 40800 53440 6 m_wbs_dat_o_1[29]
port 325 nsew signal input
rlabel metal3 s 39200 17144 40800 17264 6 m_wbs_dat_o_1[2]
port 326 nsew signal input
rlabel metal3 s 39200 54680 40800 54800 6 m_wbs_dat_o_1[30]
port 327 nsew signal input
rlabel metal3 s 39200 56040 40800 56160 6 m_wbs_dat_o_1[31]
port 328 nsew signal input
rlabel metal3 s 39200 18368 40800 18488 6 m_wbs_dat_o_1[3]
port 329 nsew signal input
rlabel metal3 s 39200 19728 40800 19848 6 m_wbs_dat_o_1[4]
port 330 nsew signal input
rlabel metal3 s 39200 21088 40800 21208 6 m_wbs_dat_o_1[5]
port 331 nsew signal input
rlabel metal3 s 39200 22448 40800 22568 6 m_wbs_dat_o_1[6]
port 332 nsew signal input
rlabel metal3 s 39200 23808 40800 23928 6 m_wbs_dat_o_1[7]
port 333 nsew signal input
rlabel metal3 s 39200 25168 40800 25288 6 m_wbs_dat_o_1[8]
port 334 nsew signal input
rlabel metal3 s 39200 26528 40800 26648 6 m_wbs_dat_o_1[9]
port 335 nsew signal input
rlabel metal3 s 39200 57400 40800 57520 6 m_wbs_dat_o_2[0]
port 336 nsew signal input
rlabel metal3 s 39200 61888 40800 62008 6 m_wbs_dat_o_2[10]
port 337 nsew signal input
rlabel metal3 s 39200 62296 40800 62416 6 m_wbs_dat_o_2[11]
port 338 nsew signal input
rlabel metal3 s 39200 62704 40800 62824 6 m_wbs_dat_o_2[12]
port 339 nsew signal input
rlabel metal3 s 39200 63248 40800 63368 6 m_wbs_dat_o_2[13]
port 340 nsew signal input
rlabel metal3 s 39200 63656 40800 63776 6 m_wbs_dat_o_2[14]
port 341 nsew signal input
rlabel metal3 s 39200 64064 40800 64184 6 m_wbs_dat_o_2[15]
port 342 nsew signal input
rlabel metal3 s 39200 64472 40800 64592 6 m_wbs_dat_o_2[16]
port 343 nsew signal input
rlabel metal3 s 39200 65016 40800 65136 6 m_wbs_dat_o_2[17]
port 344 nsew signal input
rlabel metal3 s 39200 65424 40800 65544 6 m_wbs_dat_o_2[18]
port 345 nsew signal input
rlabel metal3 s 39200 65832 40800 65952 6 m_wbs_dat_o_2[19]
port 346 nsew signal input
rlabel metal3 s 39200 57808 40800 57928 6 m_wbs_dat_o_2[1]
port 347 nsew signal input
rlabel metal3 s 39200 66376 40800 66496 6 m_wbs_dat_o_2[20]
port 348 nsew signal input
rlabel metal3 s 39200 66784 40800 66904 6 m_wbs_dat_o_2[21]
port 349 nsew signal input
rlabel metal3 s 39200 67192 40800 67312 6 m_wbs_dat_o_2[22]
port 350 nsew signal input
rlabel metal3 s 39200 67600 40800 67720 6 m_wbs_dat_o_2[23]
port 351 nsew signal input
rlabel metal3 s 39200 68144 40800 68264 6 m_wbs_dat_o_2[24]
port 352 nsew signal input
rlabel metal3 s 39200 68552 40800 68672 6 m_wbs_dat_o_2[25]
port 353 nsew signal input
rlabel metal3 s 39200 68960 40800 69080 6 m_wbs_dat_o_2[26]
port 354 nsew signal input
rlabel metal3 s 39200 69504 40800 69624 6 m_wbs_dat_o_2[27]
port 355 nsew signal input
rlabel metal3 s 39200 69912 40800 70032 6 m_wbs_dat_o_2[28]
port 356 nsew signal input
rlabel metal3 s 39200 70320 40800 70440 6 m_wbs_dat_o_2[29]
port 357 nsew signal input
rlabel metal3 s 39200 58216 40800 58336 6 m_wbs_dat_o_2[2]
port 358 nsew signal input
rlabel metal3 s 39200 70728 40800 70848 6 m_wbs_dat_o_2[30]
port 359 nsew signal input
rlabel metal3 s 39200 71272 40800 71392 6 m_wbs_dat_o_2[31]
port 360 nsew signal input
rlabel metal3 s 39200 58760 40800 58880 6 m_wbs_dat_o_2[3]
port 361 nsew signal input
rlabel metal3 s 39200 59168 40800 59288 6 m_wbs_dat_o_2[4]
port 362 nsew signal input
rlabel metal3 s 39200 59576 40800 59696 6 m_wbs_dat_o_2[5]
port 363 nsew signal input
rlabel metal3 s 39200 60120 40800 60240 6 m_wbs_dat_o_2[6]
port 364 nsew signal input
rlabel metal3 s 39200 60528 40800 60648 6 m_wbs_dat_o_2[7]
port 365 nsew signal input
rlabel metal3 s 39200 60936 40800 61056 6 m_wbs_dat_o_2[8]
port 366 nsew signal input
rlabel metal3 s 39200 61344 40800 61464 6 m_wbs_dat_o_2[9]
port 367 nsew signal input
rlabel metal3 s 39200 71680 40800 71800 6 m_wbs_dat_o_3[0]
port 368 nsew signal input
rlabel metal3 s 39200 76168 40800 76288 6 m_wbs_dat_o_3[10]
port 369 nsew signal input
rlabel metal3 s 39200 76576 40800 76696 6 m_wbs_dat_o_3[11]
port 370 nsew signal input
rlabel metal3 s 39200 77120 40800 77240 6 m_wbs_dat_o_3[12]
port 371 nsew signal input
rlabel metal3 s 39200 77528 40800 77648 6 m_wbs_dat_o_3[13]
port 372 nsew signal input
rlabel metal3 s 39200 77936 40800 78056 6 m_wbs_dat_o_3[14]
port 373 nsew signal input
rlabel metal3 s 39200 78344 40800 78464 6 m_wbs_dat_o_3[15]
port 374 nsew signal input
rlabel metal3 s 39200 78888 40800 79008 6 m_wbs_dat_o_3[16]
port 375 nsew signal input
rlabel metal3 s 39200 79296 40800 79416 6 m_wbs_dat_o_3[17]
port 376 nsew signal input
rlabel metal3 s 39200 79704 40800 79824 6 m_wbs_dat_o_3[18]
port 377 nsew signal input
rlabel metal3 s 39200 80248 40800 80368 6 m_wbs_dat_o_3[19]
port 378 nsew signal input
rlabel metal3 s 39200 72088 40800 72208 6 m_wbs_dat_o_3[1]
port 379 nsew signal input
rlabel metal3 s 39200 80656 40800 80776 6 m_wbs_dat_o_3[20]
port 380 nsew signal input
rlabel metal3 s 39200 81064 40800 81184 6 m_wbs_dat_o_3[21]
port 381 nsew signal input
rlabel metal3 s 39200 81472 40800 81592 6 m_wbs_dat_o_3[22]
port 382 nsew signal input
rlabel metal3 s 39200 82016 40800 82136 6 m_wbs_dat_o_3[23]
port 383 nsew signal input
rlabel metal3 s 39200 82424 40800 82544 6 m_wbs_dat_o_3[24]
port 384 nsew signal input
rlabel metal3 s 39200 82832 40800 82952 6 m_wbs_dat_o_3[25]
port 385 nsew signal input
rlabel metal3 s 39200 83376 40800 83496 6 m_wbs_dat_o_3[26]
port 386 nsew signal input
rlabel metal3 s 39200 83784 40800 83904 6 m_wbs_dat_o_3[27]
port 387 nsew signal input
rlabel metal3 s 39200 84192 40800 84312 6 m_wbs_dat_o_3[28]
port 388 nsew signal input
rlabel metal3 s 39200 84736 40800 84856 6 m_wbs_dat_o_3[29]
port 389 nsew signal input
rlabel metal3 s 39200 72632 40800 72752 6 m_wbs_dat_o_3[2]
port 390 nsew signal input
rlabel metal3 s 39200 85144 40800 85264 6 m_wbs_dat_o_3[30]
port 391 nsew signal input
rlabel metal3 s 39200 85552 40800 85672 6 m_wbs_dat_o_3[31]
port 392 nsew signal input
rlabel metal3 s 39200 73040 40800 73160 6 m_wbs_dat_o_3[3]
port 393 nsew signal input
rlabel metal3 s 39200 73448 40800 73568 6 m_wbs_dat_o_3[4]
port 394 nsew signal input
rlabel metal3 s 39200 73992 40800 74112 6 m_wbs_dat_o_3[5]
port 395 nsew signal input
rlabel metal3 s 39200 74400 40800 74520 6 m_wbs_dat_o_3[6]
port 396 nsew signal input
rlabel metal3 s 39200 74808 40800 74928 6 m_wbs_dat_o_3[7]
port 397 nsew signal input
rlabel metal3 s 39200 75216 40800 75336 6 m_wbs_dat_o_3[8]
port 398 nsew signal input
rlabel metal3 s 39200 75760 40800 75880 6 m_wbs_dat_o_3[9]
port 399 nsew signal input
rlabel metal3 s 39200 85960 40800 86080 6 m_wbs_dat_o_4[0]
port 400 nsew signal input
rlabel metal3 s 39200 90448 40800 90568 6 m_wbs_dat_o_4[10]
port 401 nsew signal input
rlabel metal3 s 39200 90992 40800 91112 6 m_wbs_dat_o_4[11]
port 402 nsew signal input
rlabel metal3 s 39200 91400 40800 91520 6 m_wbs_dat_o_4[12]
port 403 nsew signal input
rlabel metal3 s 39200 91808 40800 91928 6 m_wbs_dat_o_4[13]
port 404 nsew signal input
rlabel metal3 s 39200 92216 40800 92336 6 m_wbs_dat_o_4[14]
port 405 nsew signal input
rlabel metal3 s 39200 92760 40800 92880 6 m_wbs_dat_o_4[15]
port 406 nsew signal input
rlabel metal3 s 39200 93168 40800 93288 6 m_wbs_dat_o_4[16]
port 407 nsew signal input
rlabel metal3 s 39200 93576 40800 93696 6 m_wbs_dat_o_4[17]
port 408 nsew signal input
rlabel metal3 s 39200 94120 40800 94240 6 m_wbs_dat_o_4[18]
port 409 nsew signal input
rlabel metal3 s 39200 94528 40800 94648 6 m_wbs_dat_o_4[19]
port 410 nsew signal input
rlabel metal3 s 39200 86504 40800 86624 6 m_wbs_dat_o_4[1]
port 411 nsew signal input
rlabel metal3 s 39200 94936 40800 95056 6 m_wbs_dat_o_4[20]
port 412 nsew signal input
rlabel metal3 s 39200 95344 40800 95464 6 m_wbs_dat_o_4[21]
port 413 nsew signal input
rlabel metal3 s 39200 95888 40800 96008 6 m_wbs_dat_o_4[22]
port 414 nsew signal input
rlabel metal3 s 39200 96296 40800 96416 6 m_wbs_dat_o_4[23]
port 415 nsew signal input
rlabel metal3 s 39200 96704 40800 96824 6 m_wbs_dat_o_4[24]
port 416 nsew signal input
rlabel metal3 s 39200 97248 40800 97368 6 m_wbs_dat_o_4[25]
port 417 nsew signal input
rlabel metal3 s 39200 97656 40800 97776 6 m_wbs_dat_o_4[26]
port 418 nsew signal input
rlabel metal3 s 39200 98064 40800 98184 6 m_wbs_dat_o_4[27]
port 419 nsew signal input
rlabel metal3 s 39200 98608 40800 98728 6 m_wbs_dat_o_4[28]
port 420 nsew signal input
rlabel metal3 s 39200 99016 40800 99136 6 m_wbs_dat_o_4[29]
port 421 nsew signal input
rlabel metal3 s 39200 86912 40800 87032 6 m_wbs_dat_o_4[2]
port 422 nsew signal input
rlabel metal3 s 39200 99424 40800 99544 6 m_wbs_dat_o_4[30]
port 423 nsew signal input
rlabel metal3 s 39200 99832 40800 99952 6 m_wbs_dat_o_4[31]
port 424 nsew signal input
rlabel metal3 s 39200 87320 40800 87440 6 m_wbs_dat_o_4[3]
port 425 nsew signal input
rlabel metal3 s 39200 87864 40800 87984 6 m_wbs_dat_o_4[4]
port 426 nsew signal input
rlabel metal3 s 39200 88272 40800 88392 6 m_wbs_dat_o_4[5]
port 427 nsew signal input
rlabel metal3 s 39200 88680 40800 88800 6 m_wbs_dat_o_4[6]
port 428 nsew signal input
rlabel metal3 s 39200 89088 40800 89208 6 m_wbs_dat_o_4[7]
port 429 nsew signal input
rlabel metal3 s 39200 89632 40800 89752 6 m_wbs_dat_o_4[8]
port 430 nsew signal input
rlabel metal3 s 39200 90040 40800 90160 6 m_wbs_dat_o_4[9]
port 431 nsew signal input
rlabel metal3 s 39200 100376 40800 100496 6 m_wbs_dat_o_5[0]
port 432 nsew signal input
rlabel metal3 s 39200 104864 40800 104984 6 m_wbs_dat_o_5[10]
port 433 nsew signal input
rlabel metal3 s 39200 105272 40800 105392 6 m_wbs_dat_o_5[11]
port 434 nsew signal input
rlabel metal3 s 39200 105680 40800 105800 6 m_wbs_dat_o_5[12]
port 435 nsew signal input
rlabel metal3 s 39200 106088 40800 106208 6 m_wbs_dat_o_5[13]
port 436 nsew signal input
rlabel metal3 s 39200 106632 40800 106752 6 m_wbs_dat_o_5[14]
port 437 nsew signal input
rlabel metal3 s 39200 107040 40800 107160 6 m_wbs_dat_o_5[15]
port 438 nsew signal input
rlabel metal3 s 39200 107448 40800 107568 6 m_wbs_dat_o_5[16]
port 439 nsew signal input
rlabel metal3 s 39200 107992 40800 108112 6 m_wbs_dat_o_5[17]
port 440 nsew signal input
rlabel metal3 s 39200 108400 40800 108520 6 m_wbs_dat_o_5[18]
port 441 nsew signal input
rlabel metal3 s 39200 108808 40800 108928 6 m_wbs_dat_o_5[19]
port 442 nsew signal input
rlabel metal3 s 39200 100784 40800 100904 6 m_wbs_dat_o_5[1]
port 443 nsew signal input
rlabel metal3 s 39200 109352 40800 109472 6 m_wbs_dat_o_5[20]
port 444 nsew signal input
rlabel metal3 s 39200 109760 40800 109880 6 m_wbs_dat_o_5[21]
port 445 nsew signal input
rlabel metal3 s 39200 110168 40800 110288 6 m_wbs_dat_o_5[22]
port 446 nsew signal input
rlabel metal3 s 39200 110576 40800 110696 6 m_wbs_dat_o_5[23]
port 447 nsew signal input
rlabel metal3 s 39200 111120 40800 111240 6 m_wbs_dat_o_5[24]
port 448 nsew signal input
rlabel metal3 s 39200 111528 40800 111648 6 m_wbs_dat_o_5[25]
port 449 nsew signal input
rlabel metal3 s 39200 111936 40800 112056 6 m_wbs_dat_o_5[26]
port 450 nsew signal input
rlabel metal3 s 39200 112480 40800 112600 6 m_wbs_dat_o_5[27]
port 451 nsew signal input
rlabel metal3 s 39200 112888 40800 113008 6 m_wbs_dat_o_5[28]
port 452 nsew signal input
rlabel metal3 s 39200 113296 40800 113416 6 m_wbs_dat_o_5[29]
port 453 nsew signal input
rlabel metal3 s 39200 101192 40800 101312 6 m_wbs_dat_o_5[2]
port 454 nsew signal input
rlabel metal3 s 39200 113704 40800 113824 6 m_wbs_dat_o_5[30]
port 455 nsew signal input
rlabel metal3 s 39200 114248 40800 114368 6 m_wbs_dat_o_5[31]
port 456 nsew signal input
rlabel metal3 s 39200 101736 40800 101856 6 m_wbs_dat_o_5[3]
port 457 nsew signal input
rlabel metal3 s 39200 102144 40800 102264 6 m_wbs_dat_o_5[4]
port 458 nsew signal input
rlabel metal3 s 39200 102552 40800 102672 6 m_wbs_dat_o_5[5]
port 459 nsew signal input
rlabel metal3 s 39200 102960 40800 103080 6 m_wbs_dat_o_5[6]
port 460 nsew signal input
rlabel metal3 s 39200 103504 40800 103624 6 m_wbs_dat_o_5[7]
port 461 nsew signal input
rlabel metal3 s 39200 103912 40800 104032 6 m_wbs_dat_o_5[8]
port 462 nsew signal input
rlabel metal3 s 39200 104320 40800 104440 6 m_wbs_dat_o_5[9]
port 463 nsew signal input
rlabel metal3 s -800 280 800 400 4 m_wbs_dat_o_6[0]
port 464 nsew signal input
rlabel metal3 s -800 8168 800 8288 4 m_wbs_dat_o_6[10]
port 465 nsew signal input
rlabel metal3 s -800 8984 800 9104 4 m_wbs_dat_o_6[11]
port 466 nsew signal input
rlabel metal3 s -800 9800 800 9920 4 m_wbs_dat_o_6[12]
port 467 nsew signal input
rlabel metal3 s -800 10616 800 10736 4 m_wbs_dat_o_6[13]
port 468 nsew signal input
rlabel metal3 s -800 11432 800 11552 4 m_wbs_dat_o_6[14]
port 469 nsew signal input
rlabel metal3 s -800 12248 800 12368 4 m_wbs_dat_o_6[15]
port 470 nsew signal input
rlabel metal3 s -800 13064 800 13184 4 m_wbs_dat_o_6[16]
port 471 nsew signal input
rlabel metal3 s -800 13744 800 13864 4 m_wbs_dat_o_6[17]
port 472 nsew signal input
rlabel metal3 s -800 14560 800 14680 4 m_wbs_dat_o_6[18]
port 473 nsew signal input
rlabel metal3 s -800 15376 800 15496 4 m_wbs_dat_o_6[19]
port 474 nsew signal input
rlabel metal3 s -800 960 800 1080 4 m_wbs_dat_o_6[1]
port 475 nsew signal input
rlabel metal3 s -800 16192 800 16312 4 m_wbs_dat_o_6[20]
port 476 nsew signal input
rlabel metal3 s -800 17008 800 17128 4 m_wbs_dat_o_6[21]
port 477 nsew signal input
rlabel metal3 s -800 17824 800 17944 4 m_wbs_dat_o_6[22]
port 478 nsew signal input
rlabel metal3 s -800 18640 800 18760 4 m_wbs_dat_o_6[23]
port 479 nsew signal input
rlabel metal3 s -800 19456 800 19576 4 m_wbs_dat_o_6[24]
port 480 nsew signal input
rlabel metal3 s -800 20272 800 20392 4 m_wbs_dat_o_6[25]
port 481 nsew signal input
rlabel metal3 s -800 20952 800 21072 4 m_wbs_dat_o_6[26]
port 482 nsew signal input
rlabel metal3 s -800 21768 800 21888 4 m_wbs_dat_o_6[27]
port 483 nsew signal input
rlabel metal3 s -800 22584 800 22704 4 m_wbs_dat_o_6[28]
port 484 nsew signal input
rlabel metal3 s -800 23400 800 23520 4 m_wbs_dat_o_6[29]
port 485 nsew signal input
rlabel metal3 s -800 1776 800 1896 4 m_wbs_dat_o_6[2]
port 486 nsew signal input
rlabel metal3 s -800 24216 800 24336 4 m_wbs_dat_o_6[30]
port 487 nsew signal input
rlabel metal3 s -800 25032 800 25152 4 m_wbs_dat_o_6[31]
port 488 nsew signal input
rlabel metal3 s -800 2592 800 2712 4 m_wbs_dat_o_6[3]
port 489 nsew signal input
rlabel metal3 s -800 3408 800 3528 4 m_wbs_dat_o_6[4]
port 490 nsew signal input
rlabel metal3 s -800 4224 800 4344 4 m_wbs_dat_o_6[5]
port 491 nsew signal input
rlabel metal3 s -800 5040 800 5160 4 m_wbs_dat_o_6[6]
port 492 nsew signal input
rlabel metal3 s -800 5856 800 5976 4 m_wbs_dat_o_6[7]
port 493 nsew signal input
rlabel metal3 s -800 6672 800 6792 4 m_wbs_dat_o_6[8]
port 494 nsew signal input
rlabel metal3 s -800 7352 800 7472 4 m_wbs_dat_o_6[9]
port 495 nsew signal input
rlabel metal3 s -800 25848 800 25968 4 m_wbs_dat_o_7[0]
port 496 nsew signal input
rlabel metal3 s -800 33736 800 33856 4 m_wbs_dat_o_7[10]
port 497 nsew signal input
rlabel metal3 s -800 34552 800 34672 4 m_wbs_dat_o_7[11]
port 498 nsew signal input
rlabel metal3 s -800 35368 800 35488 4 m_wbs_dat_o_7[12]
port 499 nsew signal input
rlabel metal3 s -800 36184 800 36304 4 m_wbs_dat_o_7[13]
port 500 nsew signal input
rlabel metal3 s -800 37000 800 37120 4 m_wbs_dat_o_7[14]
port 501 nsew signal input
rlabel metal3 s -800 37816 800 37936 4 m_wbs_dat_o_7[15]
port 502 nsew signal input
rlabel metal3 s -800 38632 800 38752 4 m_wbs_dat_o_7[16]
port 503 nsew signal input
rlabel metal3 s -800 39448 800 39568 4 m_wbs_dat_o_7[17]
port 504 nsew signal input
rlabel metal3 s -800 40264 800 40384 4 m_wbs_dat_o_7[18]
port 505 nsew signal input
rlabel metal3 s -800 40944 800 41064 4 m_wbs_dat_o_7[19]
port 506 nsew signal input
rlabel metal3 s -800 26664 800 26784 4 m_wbs_dat_o_7[1]
port 507 nsew signal input
rlabel metal3 s -800 41760 800 41880 4 m_wbs_dat_o_7[20]
port 508 nsew signal input
rlabel metal3 s -800 42576 800 42696 4 m_wbs_dat_o_7[21]
port 509 nsew signal input
rlabel metal3 s -800 43392 800 43512 4 m_wbs_dat_o_7[22]
port 510 nsew signal input
rlabel metal3 s -800 44208 800 44328 4 m_wbs_dat_o_7[23]
port 511 nsew signal input
rlabel metal3 s -800 45024 800 45144 4 m_wbs_dat_o_7[24]
port 512 nsew signal input
rlabel metal3 s -800 45840 800 45960 4 m_wbs_dat_o_7[25]
port 513 nsew signal input
rlabel metal3 s -800 46656 800 46776 4 m_wbs_dat_o_7[26]
port 514 nsew signal input
rlabel metal3 s -800 47336 800 47456 4 m_wbs_dat_o_7[27]
port 515 nsew signal input
rlabel metal3 s -800 48152 800 48272 4 m_wbs_dat_o_7[28]
port 516 nsew signal input
rlabel metal3 s -800 48968 800 49088 4 m_wbs_dat_o_7[29]
port 517 nsew signal input
rlabel metal3 s -800 27344 800 27464 4 m_wbs_dat_o_7[2]
port 518 nsew signal input
rlabel metal3 s -800 49784 800 49904 4 m_wbs_dat_o_7[30]
port 519 nsew signal input
rlabel metal3 s -800 50600 800 50720 4 m_wbs_dat_o_7[31]
port 520 nsew signal input
rlabel metal3 s -800 28160 800 28280 4 m_wbs_dat_o_7[3]
port 521 nsew signal input
rlabel metal3 s -800 28976 800 29096 4 m_wbs_dat_o_7[4]
port 522 nsew signal input
rlabel metal3 s -800 29792 800 29912 4 m_wbs_dat_o_7[5]
port 523 nsew signal input
rlabel metal3 s -800 30608 800 30728 4 m_wbs_dat_o_7[6]
port 524 nsew signal input
rlabel metal3 s -800 31424 800 31544 4 m_wbs_dat_o_7[7]
port 525 nsew signal input
rlabel metal3 s -800 32240 800 32360 4 m_wbs_dat_o_7[8]
port 526 nsew signal input
rlabel metal3 s -800 33056 800 33176 4 m_wbs_dat_o_7[9]
port 527 nsew signal input
rlabel metal3 s -800 51416 800 51536 4 m_wbs_dat_o_8[0]
port 528 nsew signal input
rlabel metal3 s -800 59440 800 59560 4 m_wbs_dat_o_8[10]
port 529 nsew signal input
rlabel metal3 s -800 60256 800 60376 4 m_wbs_dat_o_8[11]
port 530 nsew signal input
rlabel metal3 s -800 60936 800 61056 4 m_wbs_dat_o_8[12]
port 531 nsew signal input
rlabel metal3 s -800 61752 800 61872 4 m_wbs_dat_o_8[13]
port 532 nsew signal input
rlabel metal3 s -800 62568 800 62688 4 m_wbs_dat_o_8[14]
port 533 nsew signal input
rlabel metal3 s -800 63384 800 63504 4 m_wbs_dat_o_8[15]
port 534 nsew signal input
rlabel metal3 s -800 64200 800 64320 4 m_wbs_dat_o_8[16]
port 535 nsew signal input
rlabel metal3 s -800 65016 800 65136 4 m_wbs_dat_o_8[17]
port 536 nsew signal input
rlabel metal3 s -800 65832 800 65952 4 m_wbs_dat_o_8[18]
port 537 nsew signal input
rlabel metal3 s -800 66648 800 66768 4 m_wbs_dat_o_8[19]
port 538 nsew signal input
rlabel metal3 s -800 52232 800 52352 4 m_wbs_dat_o_8[1]
port 539 nsew signal input
rlabel metal3 s -800 67328 800 67448 4 m_wbs_dat_o_8[20]
port 540 nsew signal input
rlabel metal3 s -800 68144 800 68264 4 m_wbs_dat_o_8[21]
port 541 nsew signal input
rlabel metal3 s -800 68960 800 69080 4 m_wbs_dat_o_8[22]
port 542 nsew signal input
rlabel metal3 s -800 69776 800 69896 4 m_wbs_dat_o_8[23]
port 543 nsew signal input
rlabel metal3 s -800 70592 800 70712 4 m_wbs_dat_o_8[24]
port 544 nsew signal input
rlabel metal3 s -800 71408 800 71528 4 m_wbs_dat_o_8[25]
port 545 nsew signal input
rlabel metal3 s -800 72224 800 72344 4 m_wbs_dat_o_8[26]
port 546 nsew signal input
rlabel metal3 s -800 73040 800 73160 4 m_wbs_dat_o_8[27]
port 547 nsew signal input
rlabel metal3 s -800 73720 800 73840 4 m_wbs_dat_o_8[28]
port 548 nsew signal input
rlabel metal3 s -800 74536 800 74656 4 m_wbs_dat_o_8[29]
port 549 nsew signal input
rlabel metal3 s -800 53048 800 53168 4 m_wbs_dat_o_8[2]
port 550 nsew signal input
rlabel metal3 s -800 75352 800 75472 4 m_wbs_dat_o_8[30]
port 551 nsew signal input
rlabel metal3 s -800 76168 800 76288 4 m_wbs_dat_o_8[31]
port 552 nsew signal input
rlabel metal3 s -800 53728 800 53848 4 m_wbs_dat_o_8[3]
port 553 nsew signal input
rlabel metal3 s -800 54544 800 54664 4 m_wbs_dat_o_8[4]
port 554 nsew signal input
rlabel metal3 s -800 55360 800 55480 4 m_wbs_dat_o_8[5]
port 555 nsew signal input
rlabel metal3 s -800 56176 800 56296 4 m_wbs_dat_o_8[6]
port 556 nsew signal input
rlabel metal3 s -800 56992 800 57112 4 m_wbs_dat_o_8[7]
port 557 nsew signal input
rlabel metal3 s -800 57808 800 57928 4 m_wbs_dat_o_8[8]
port 558 nsew signal input
rlabel metal3 s -800 58624 800 58744 4 m_wbs_dat_o_8[9]
port 559 nsew signal input
rlabel metal3 s -800 76984 800 77104 4 m_wbs_dat_o_9[0]
port 560 nsew signal input
rlabel metal3 s -800 85008 800 85128 4 m_wbs_dat_o_9[10]
port 561 nsew signal input
rlabel metal3 s -800 85824 800 85944 4 m_wbs_dat_o_9[11]
port 562 nsew signal input
rlabel metal3 s -800 86640 800 86760 4 m_wbs_dat_o_9[12]
port 563 nsew signal input
rlabel metal3 s -800 87320 800 87440 4 m_wbs_dat_o_9[13]
port 564 nsew signal input
rlabel metal3 s -800 88136 800 88256 4 m_wbs_dat_o_9[14]
port 565 nsew signal input
rlabel metal3 s -800 88952 800 89072 4 m_wbs_dat_o_9[15]
port 566 nsew signal input
rlabel metal3 s -800 89768 800 89888 4 m_wbs_dat_o_9[16]
port 567 nsew signal input
rlabel metal3 s -800 90584 800 90704 4 m_wbs_dat_o_9[17]
port 568 nsew signal input
rlabel metal3 s -800 91400 800 91520 4 m_wbs_dat_o_9[18]
port 569 nsew signal input
rlabel metal3 s -800 92216 800 92336 4 m_wbs_dat_o_9[19]
port 570 nsew signal input
rlabel metal3 s -800 77800 800 77920 4 m_wbs_dat_o_9[1]
port 571 nsew signal input
rlabel metal3 s -800 93032 800 93152 4 m_wbs_dat_o_9[20]
port 572 nsew signal input
rlabel metal3 s -800 93712 800 93832 4 m_wbs_dat_o_9[21]
port 573 nsew signal input
rlabel metal3 s -800 94528 800 94648 4 m_wbs_dat_o_9[22]
port 574 nsew signal input
rlabel metal3 s -800 95344 800 95464 4 m_wbs_dat_o_9[23]
port 575 nsew signal input
rlabel metal3 s -800 96160 800 96280 4 m_wbs_dat_o_9[24]
port 576 nsew signal input
rlabel metal3 s -800 96976 800 97096 4 m_wbs_dat_o_9[25]
port 577 nsew signal input
rlabel metal3 s -800 97792 800 97912 4 m_wbs_dat_o_9[26]
port 578 nsew signal input
rlabel metal3 s -800 98608 800 98728 4 m_wbs_dat_o_9[27]
port 579 nsew signal input
rlabel metal3 s -800 99424 800 99544 4 m_wbs_dat_o_9[28]
port 580 nsew signal input
rlabel metal3 s -800 100240 800 100360 4 m_wbs_dat_o_9[29]
port 581 nsew signal input
rlabel metal3 s -800 78616 800 78736 4 m_wbs_dat_o_9[2]
port 582 nsew signal input
rlabel metal3 s -800 100920 800 101040 4 m_wbs_dat_o_9[30]
port 583 nsew signal input
rlabel metal3 s -800 101736 800 101856 4 m_wbs_dat_o_9[31]
port 584 nsew signal input
rlabel metal3 s -800 79432 800 79552 4 m_wbs_dat_o_9[3]
port 585 nsew signal input
rlabel metal3 s -800 80248 800 80368 4 m_wbs_dat_o_9[4]
port 586 nsew signal input
rlabel metal3 s -800 80928 800 81048 4 m_wbs_dat_o_9[5]
port 587 nsew signal input
rlabel metal3 s -800 81744 800 81864 4 m_wbs_dat_o_9[6]
port 588 nsew signal input
rlabel metal3 s -800 82560 800 82680 4 m_wbs_dat_o_9[7]
port 589 nsew signal input
rlabel metal3 s -800 83376 800 83496 4 m_wbs_dat_o_9[8]
port 590 nsew signal input
rlabel metal3 s -800 84192 800 84312 4 m_wbs_dat_o_9[9]
port 591 nsew signal input
rlabel metal3 s -800 102552 800 102672 4 m_wbs_we_i
port 592 nsew signal output
rlabel metal2 s 28262 119200 28318 120800 6 mt_QEI_ChA_0
port 593 nsew signal output
rlabel metal2 s 28538 119200 28594 120800 6 mt_QEI_ChA_1
port 594 nsew signal output
rlabel metal2 s 28722 119200 28778 120800 6 mt_QEI_ChA_2
port 595 nsew signal output
rlabel metal2 s 28998 119200 29054 120800 6 mt_QEI_ChA_3
port 596 nsew signal output
rlabel metal2 s 29182 119200 29238 120800 6 mt_QEI_ChB_0
port 597 nsew signal output
rlabel metal2 s 29458 119200 29514 120800 6 mt_QEI_ChB_1
port 598 nsew signal output
rlabel metal2 s 29642 119200 29698 120800 6 mt_QEI_ChB_2
port 599 nsew signal output
rlabel metal2 s 29918 119200 29974 120800 6 mt_QEI_ChB_3
port 600 nsew signal output
rlabel metal2 s 30102 119200 30158 120800 6 mt_pwm_h_0
port 601 nsew signal input
rlabel metal2 s 30378 119200 30434 120800 6 mt_pwm_h_1
port 602 nsew signal input
rlabel metal2 s 30562 119200 30618 120800 6 mt_pwm_h_2
port 603 nsew signal input
rlabel metal2 s 30838 119200 30894 120800 6 mt_pwm_h_3
port 604 nsew signal input
rlabel metal2 s 31022 119200 31078 120800 6 mt_pwm_l_0
port 605 nsew signal input
rlabel metal2 s 31298 119200 31354 120800 6 mt_pwm_l_1
port 606 nsew signal input
rlabel metal2 s 31482 119200 31538 120800 6 mt_pwm_l_2
port 607 nsew signal input
rlabel metal2 s 31758 119200 31814 120800 6 mt_pwm_l_3
port 608 nsew signal input
rlabel metal2 s 110 -800 166 800 8 wb_clk_i
port 609 nsew signal input
rlabel metal2 s 386 -800 442 800 8 wb_rst_i
port 610 nsew signal input
rlabel metal2 s 1674 -800 1730 800 8 wbs_ack_o
port 611 nsew signal output
rlabel metal2 s 2962 -800 3018 800 8 wbs_adr_i[0]
port 612 nsew signal input
rlabel metal2 s 14094 -800 14150 800 8 wbs_adr_i[10]
port 613 nsew signal input
rlabel metal2 s 15014 -800 15070 800 8 wbs_adr_i[11]
port 614 nsew signal input
rlabel metal2 s 16026 -800 16082 800 8 wbs_adr_i[12]
port 615 nsew signal input
rlabel metal2 s 16946 -800 17002 800 8 wbs_adr_i[13]
port 616 nsew signal input
rlabel metal2 s 17958 -800 18014 800 8 wbs_adr_i[14]
port 617 nsew signal input
rlabel metal2 s 18970 -800 19026 800 8 wbs_adr_i[15]
port 618 nsew signal input
rlabel metal2 s 19890 -800 19946 800 8 wbs_adr_i[16]
port 619 nsew signal input
rlabel metal2 s 20902 -800 20958 800 8 wbs_adr_i[17]
port 620 nsew signal input
rlabel metal2 s 21822 -800 21878 800 8 wbs_adr_i[18]
port 621 nsew signal input
rlabel metal2 s 22834 -800 22890 800 8 wbs_adr_i[19]
port 622 nsew signal input
rlabel metal2 s 4250 -800 4306 800 8 wbs_adr_i[1]
port 623 nsew signal input
rlabel metal2 s 23846 -800 23902 800 8 wbs_adr_i[20]
port 624 nsew signal input
rlabel metal2 s 24766 -800 24822 800 8 wbs_adr_i[21]
port 625 nsew signal input
rlabel metal2 s 25778 -800 25834 800 8 wbs_adr_i[22]
port 626 nsew signal input
rlabel metal2 s 26790 -800 26846 800 8 wbs_adr_i[23]
port 627 nsew signal input
rlabel metal2 s 27710 -800 27766 800 8 wbs_adr_i[24]
port 628 nsew signal input
rlabel metal2 s 28722 -800 28778 800 8 wbs_adr_i[25]
port 629 nsew signal input
rlabel metal2 s 29642 -800 29698 800 8 wbs_adr_i[26]
port 630 nsew signal input
rlabel metal2 s 30654 -800 30710 800 8 wbs_adr_i[27]
port 631 nsew signal input
rlabel metal2 s 31666 -800 31722 800 8 wbs_adr_i[28]
port 632 nsew signal input
rlabel metal2 s 32586 -800 32642 800 8 wbs_adr_i[29]
port 633 nsew signal input
rlabel metal2 s 5630 -800 5686 800 8 wbs_adr_i[2]
port 634 nsew signal input
rlabel metal2 s 33598 -800 33654 800 8 wbs_adr_i[30]
port 635 nsew signal input
rlabel metal2 s 34518 -800 34574 800 8 wbs_adr_i[31]
port 636 nsew signal input
rlabel metal2 s 6918 -800 6974 800 8 wbs_adr_i[3]
port 637 nsew signal input
rlabel metal2 s 8206 -800 8262 800 8 wbs_adr_i[4]
port 638 nsew signal input
rlabel metal2 s 9218 -800 9274 800 8 wbs_adr_i[5]
port 639 nsew signal input
rlabel metal2 s 10138 -800 10194 800 8 wbs_adr_i[6]
port 640 nsew signal input
rlabel metal2 s 11150 -800 11206 800 8 wbs_adr_i[7]
port 641 nsew signal input
rlabel metal2 s 12070 -800 12126 800 8 wbs_adr_i[8]
port 642 nsew signal input
rlabel metal2 s 13082 -800 13138 800 8 wbs_adr_i[9]
port 643 nsew signal input
rlabel metal2 s 2042 -800 2098 800 8 wbs_cyc_i
port 644 nsew signal input
rlabel metal2 s 3330 -800 3386 800 8 wbs_dat_i[0]
port 645 nsew signal input
rlabel metal2 s 14370 -800 14426 800 8 wbs_dat_i[10]
port 646 nsew signal input
rlabel metal2 s 15382 -800 15438 800 8 wbs_dat_i[11]
port 647 nsew signal input
rlabel metal2 s 16302 -800 16358 800 8 wbs_dat_i[12]
port 648 nsew signal input
rlabel metal2 s 17314 -800 17370 800 8 wbs_dat_i[13]
port 649 nsew signal input
rlabel metal2 s 18326 -800 18382 800 8 wbs_dat_i[14]
port 650 nsew signal input
rlabel metal2 s 19246 -800 19302 800 8 wbs_dat_i[15]
port 651 nsew signal input
rlabel metal2 s 20258 -800 20314 800 8 wbs_dat_i[16]
port 652 nsew signal input
rlabel metal2 s 21178 -800 21234 800 8 wbs_dat_i[17]
port 653 nsew signal input
rlabel metal2 s 22190 -800 22246 800 8 wbs_dat_i[18]
port 654 nsew signal input
rlabel metal2 s 23202 -800 23258 800 8 wbs_dat_i[19]
port 655 nsew signal input
rlabel metal2 s 4618 -800 4674 800 8 wbs_dat_i[1]
port 656 nsew signal input
rlabel metal2 s 24122 -800 24178 800 8 wbs_dat_i[20]
port 657 nsew signal input
rlabel metal2 s 25134 -800 25190 800 8 wbs_dat_i[21]
port 658 nsew signal input
rlabel metal2 s 26054 -800 26110 800 8 wbs_dat_i[22]
port 659 nsew signal input
rlabel metal2 s 27066 -800 27122 800 8 wbs_dat_i[23]
port 660 nsew signal input
rlabel metal2 s 28078 -800 28134 800 8 wbs_dat_i[24]
port 661 nsew signal input
rlabel metal2 s 28998 -800 29054 800 8 wbs_dat_i[25]
port 662 nsew signal input
rlabel metal2 s 30010 -800 30066 800 8 wbs_dat_i[26]
port 663 nsew signal input
rlabel metal2 s 30930 -800 30986 800 8 wbs_dat_i[27]
port 664 nsew signal input
rlabel metal2 s 31942 -800 31998 800 8 wbs_dat_i[28]
port 665 nsew signal input
rlabel metal2 s 32954 -800 33010 800 8 wbs_dat_i[29]
port 666 nsew signal input
rlabel metal2 s 5906 -800 5962 800 8 wbs_dat_i[2]
port 667 nsew signal input
rlabel metal2 s 33874 -800 33930 800 8 wbs_dat_i[30]
port 668 nsew signal input
rlabel metal2 s 34886 -800 34942 800 8 wbs_dat_i[31]
port 669 nsew signal input
rlabel metal2 s 7194 -800 7250 800 8 wbs_dat_i[3]
port 670 nsew signal input
rlabel metal2 s 8482 -800 8538 800 8 wbs_dat_i[4]
port 671 nsew signal input
rlabel metal2 s 9494 -800 9550 800 8 wbs_dat_i[5]
port 672 nsew signal input
rlabel metal2 s 10506 -800 10562 800 8 wbs_dat_i[6]
port 673 nsew signal input
rlabel metal2 s 11426 -800 11482 800 8 wbs_dat_i[7]
port 674 nsew signal input
rlabel metal2 s 12438 -800 12494 800 8 wbs_dat_i[8]
port 675 nsew signal input
rlabel metal2 s 13450 -800 13506 800 8 wbs_dat_i[9]
port 676 nsew signal input
rlabel metal2 s 3606 -800 3662 800 8 wbs_dat_o[0]
port 677 nsew signal output
rlabel metal2 s 14738 -800 14794 800 8 wbs_dat_o[10]
port 678 nsew signal output
rlabel metal2 s 15658 -800 15714 800 8 wbs_dat_o[11]
port 679 nsew signal output
rlabel metal2 s 16670 -800 16726 800 8 wbs_dat_o[12]
port 680 nsew signal output
rlabel metal2 s 17590 -800 17646 800 8 wbs_dat_o[13]
port 681 nsew signal output
rlabel metal2 s 18602 -800 18658 800 8 wbs_dat_o[14]
port 682 nsew signal output
rlabel metal2 s 19614 -800 19670 800 8 wbs_dat_o[15]
port 683 nsew signal output
rlabel metal2 s 20534 -800 20590 800 8 wbs_dat_o[16]
port 684 nsew signal output
rlabel metal2 s 21546 -800 21602 800 8 wbs_dat_o[17]
port 685 nsew signal output
rlabel metal2 s 22558 -800 22614 800 8 wbs_dat_o[18]
port 686 nsew signal output
rlabel metal2 s 23478 -800 23534 800 8 wbs_dat_o[19]
port 687 nsew signal output
rlabel metal2 s 4986 -800 5042 800 8 wbs_dat_o[1]
port 688 nsew signal output
rlabel metal2 s 24490 -800 24546 800 8 wbs_dat_o[20]
port 689 nsew signal output
rlabel metal2 s 25410 -800 25466 800 8 wbs_dat_o[21]
port 690 nsew signal output
rlabel metal2 s 26422 -800 26478 800 8 wbs_dat_o[22]
port 691 nsew signal output
rlabel metal2 s 27434 -800 27490 800 8 wbs_dat_o[23]
port 692 nsew signal output
rlabel metal2 s 28354 -800 28410 800 8 wbs_dat_o[24]
port 693 nsew signal output
rlabel metal2 s 29366 -800 29422 800 8 wbs_dat_o[25]
port 694 nsew signal output
rlabel metal2 s 30286 -800 30342 800 8 wbs_dat_o[26]
port 695 nsew signal output
rlabel metal2 s 31298 -800 31354 800 8 wbs_dat_o[27]
port 696 nsew signal output
rlabel metal2 s 32310 -800 32366 800 8 wbs_dat_o[28]
port 697 nsew signal output
rlabel metal2 s 33230 -800 33286 800 8 wbs_dat_o[29]
port 698 nsew signal output
rlabel metal2 s 6274 -800 6330 800 8 wbs_dat_o[2]
port 699 nsew signal output
rlabel metal2 s 34242 -800 34298 800 8 wbs_dat_o[30]
port 700 nsew signal output
rlabel metal2 s 35162 -800 35218 800 8 wbs_dat_o[31]
port 701 nsew signal output
rlabel metal2 s 7562 -800 7618 800 8 wbs_dat_o[3]
port 702 nsew signal output
rlabel metal2 s 8850 -800 8906 800 8 wbs_dat_o[4]
port 703 nsew signal output
rlabel metal2 s 9862 -800 9918 800 8 wbs_dat_o[5]
port 704 nsew signal output
rlabel metal2 s 10782 -800 10838 800 8 wbs_dat_o[6]
port 705 nsew signal output
rlabel metal2 s 11794 -800 11850 800 8 wbs_dat_o[7]
port 706 nsew signal output
rlabel metal2 s 12714 -800 12770 800 8 wbs_dat_o[8]
port 707 nsew signal output
rlabel metal2 s 13726 -800 13782 800 8 wbs_dat_o[9]
port 708 nsew signal output
rlabel metal2 s 3974 -800 4030 800 8 wbs_sel_i[0]
port 709 nsew signal input
rlabel metal2 s 5262 -800 5318 800 8 wbs_sel_i[1]
port 710 nsew signal input
rlabel metal2 s 6550 -800 6606 800 8 wbs_sel_i[2]
port 711 nsew signal input
rlabel metal2 s 7838 -800 7894 800 8 wbs_sel_i[3]
port 712 nsew signal input
rlabel metal2 s 2318 -800 2374 800 8 wbs_stb_i
port 713 nsew signal input
rlabel metal2 s 2686 -800 2742 800 8 wbs_we_i
port 714 nsew signal input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 715 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 716 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 717 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 40000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/wb_local/runs/wb_local/results/magic/wb_local.gds
string GDS_END 3948798
string GDS_START 325112
<< end >>

