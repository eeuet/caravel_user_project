* NGSPICE file created from motor_top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

.subckt motor_top clock io_QEI_ChA io_QEI_ChB io_irq io_pwm_h io_pwm_l io_wb_ack_o
+ io_wb_adr_i[0] io_wb_adr_i[10] io_wb_adr_i[11] io_wb_adr_i[1] io_wb_adr_i[2] io_wb_adr_i[3]
+ io_wb_adr_i[4] io_wb_adr_i[5] io_wb_adr_i[6] io_wb_adr_i[7] io_wb_adr_i[8] io_wb_adr_i[9]
+ io_wb_cs_i io_wb_dat_i[0] io_wb_dat_i[10] io_wb_dat_i[11] io_wb_dat_i[12] io_wb_dat_i[13]
+ io_wb_dat_i[14] io_wb_dat_i[15] io_wb_dat_i[16] io_wb_dat_i[17] io_wb_dat_i[18]
+ io_wb_dat_i[19] io_wb_dat_i[1] io_wb_dat_i[20] io_wb_dat_i[21] io_wb_dat_i[22] io_wb_dat_i[23]
+ io_wb_dat_i[24] io_wb_dat_i[25] io_wb_dat_i[26] io_wb_dat_i[27] io_wb_dat_i[28]
+ io_wb_dat_i[29] io_wb_dat_i[2] io_wb_dat_i[30] io_wb_dat_i[31] io_wb_dat_i[3] io_wb_dat_i[4]
+ io_wb_dat_i[5] io_wb_dat_i[6] io_wb_dat_i[7] io_wb_dat_i[8] io_wb_dat_i[9] io_wb_dat_o[0]
+ io_wb_dat_o[10] io_wb_dat_o[11] io_wb_dat_o[12] io_wb_dat_o[13] io_wb_dat_o[14]
+ io_wb_dat_o[15] io_wb_dat_o[16] io_wb_dat_o[17] io_wb_dat_o[18] io_wb_dat_o[19]
+ io_wb_dat_o[1] io_wb_dat_o[20] io_wb_dat_o[21] io_wb_dat_o[22] io_wb_dat_o[23] io_wb_dat_o[24]
+ io_wb_dat_o[25] io_wb_dat_o[26] io_wb_dat_o[27] io_wb_dat_o[28] io_wb_dat_o[29]
+ io_wb_dat_o[2] io_wb_dat_o[30] io_wb_dat_o[31] io_wb_dat_o[3] io_wb_dat_o[4] io_wb_dat_o[5]
+ io_wb_dat_o[6] io_wb_dat_o[7] io_wb_dat_o[8] io_wb_dat_o[9] io_wb_we_i reset vccd1
+ vssd1
XFILLER_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7963_ _7991_/A vssd1 vssd1 vccd1 vccd1 _7987_/B sky130_fd_sc_hd__buf_1
X_9702_ _9819_/CLK _9702_/D vssd1 vssd1 vccd1 vccd1 _9702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6914_ _6907_/X _6908_/X _6907_/X _6908_/X vssd1 vssd1 vccd1 vccd1 _6914_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7894_ _7892_/A _7892_/B _7790_/X _7893_/Y vssd1 vssd1 vccd1 vccd1 _7894_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9633_ _9708_/CLK _9633_/D vssd1 vssd1 vccd1 vccd1 _9633_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6845_ _6829_/A _6835_/A _6829_/Y vssd1 vssd1 vccd1 vccd1 _6845_/X sky130_fd_sc_hd__a21o_1
XFILLER_195_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9564_ _9761_/CLK _9564_/D vssd1 vssd1 vccd1 vccd1 _9564_/Q sky130_fd_sc_hd__dfxtp_1
X_6776_ _6766_/C _6775_/A _6765_/A _6775_/Y vssd1 vssd1 vccd1 vccd1 _6776_/X sky130_fd_sc_hd__a22o_1
X_8515_ _8481_/X _8514_/X _8481_/X _8514_/X vssd1 vssd1 vccd1 vccd1 _8515_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_148_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5727_ _6576_/A _9660_/Q _5725_/A _5726_/Y vssd1 vssd1 vccd1 vccd1 _5727_/X sky130_fd_sc_hd__a22o_1
X_9495_ _7941_/X _5997_/B _9504_/S vssd1 vssd1 vccd1 vccd1 _9495_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8446_ _8446_/A _8446_/B vssd1 vssd1 vccd1 vccd1 _8467_/A sky130_fd_sc_hd__or2_1
XFILLER_136_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5658_ _5689_/A vssd1 vssd1 vccd1 vccd1 _5658_/X sky130_fd_sc_hd__clkbuf_2
X_8377_ _8377_/A _8377_/B vssd1 vssd1 vccd1 vccd1 _9561_/D sky130_fd_sc_hd__and2_1
XFILLER_184_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5589_ _9708_/Q vssd1 vssd1 vccd1 vccd1 _7646_/A sky130_fd_sc_hd__inv_2
XFILLER_2_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7328_ _7385_/B vssd1 vssd1 vccd1 vccd1 _7400_/B sky130_fd_sc_hd__buf_1
XFILLER_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7259_ _7259_/A _7259_/B vssd1 vssd1 vccd1 vccd1 _7260_/B sky130_fd_sc_hd__or2_2
XFILLER_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4960_ _9847_/Q vssd1 vssd1 vccd1 vccd1 _4960_/X sky130_fd_sc_hd__buf_2
X_4891_ _9732_/Q _4865_/X _9880_/Q _4866_/X _4887_/X vssd1 vssd1 vccd1 vccd1 _9880_/D
+ sky130_fd_sc_hd__a221o_1
X_6630_ _6660_/A _6969_/B _6981_/A _9462_/X vssd1 vssd1 vccd1 vccd1 _6630_/X sky130_fd_sc_hd__or4_4
XFILLER_149_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6561_ _6561_/A vssd1 vssd1 vccd1 vccd1 _6561_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8300_ _4765_/A _8301_/B _4770_/X _8198_/X vssd1 vssd1 vccd1 vccd1 _8302_/B sky130_fd_sc_hd__o22a_1
Xrepeater93 _9306_/S vssd1 vssd1 vccd1 vccd1 _9334_/S sky130_fd_sc_hd__buf_4
XFILLER_164_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5512_ _7160_/A _7389_/B _6867_/C _6642_/A vssd1 vssd1 vccd1 vccd1 _5513_/A sky130_fd_sc_hd__o22a_1
XFILLER_118_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6492_ _6432_/Y _6460_/Y _6466_/Y _6491_/X _6465_/D vssd1 vssd1 vccd1 vccd1 _6492_/X
+ sky130_fd_sc_hd__o221a_1
X_9280_ _9763_/Q _9279_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9280_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8231_ _8231_/A _8231_/B vssd1 vssd1 vccd1 vccd1 _8232_/B sky130_fd_sc_hd__or2_1
X_5443_ _6796_/C _5442_/B _5442_/Y vssd1 vssd1 vccd1 vccd1 _7321_/D sky130_fd_sc_hd__a21oi_4
XFILLER_145_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8162_ _4802_/A _8105_/Y _4798_/A _8104_/X _8161_/X vssd1 vssd1 vccd1 vccd1 _8162_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5374_ _5374_/A vssd1 vssd1 vccd1 vccd1 _9724_/D sky130_fd_sc_hd__inv_2
X_7113_ _7334_/A vssd1 vssd1 vccd1 vccd1 _7311_/A sky130_fd_sc_hd__clkbuf_2
X_8093_ _8093_/A vssd1 vssd1 vccd1 vccd1 _8093_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7044_ _7028_/X _7030_/X _7028_/X _7030_/X vssd1 vssd1 vccd1 vccd1 _7061_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8995_ _9528_/Q _5035_/A _9445_/S vssd1 vssd1 vccd1 vccd1 _8995_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7946_ _8875_/A vssd1 vssd1 vccd1 vccd1 _8959_/A sky130_fd_sc_hd__buf_2
XFILLER_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7877_ _7877_/A _7877_/B vssd1 vssd1 vccd1 vccd1 _7882_/B sky130_fd_sc_hd__or2_2
XFILLER_42_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9616_ _9656_/CLK _9616_/D vssd1 vssd1 vccd1 vccd1 _9616_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6828_ _6813_/A _6823_/Y _6820_/X _6824_/X vssd1 vssd1 vccd1 vccd1 _6835_/A sky130_fd_sc_hd__o22ai_4
XFILLER_195_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9547_ _9916_/CLK _9547_/D vssd1 vssd1 vccd1 vccd1 _9547_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6759_ _6759_/A _6759_/B vssd1 vssd1 vccd1 vccd1 _6759_/X sky130_fd_sc_hd__or2_1
X_9478_ _6316_/B _7906_/A _9480_/S vssd1 vssd1 vccd1 vccd1 _9478_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8429_ _8436_/C _8427_/X _8440_/A vssd1 vssd1 vccd1 vccd1 _8429_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_151_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5090_ _9834_/Q vssd1 vssd1 vccd1 vccd1 _5090_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8780_ _8778_/X _8805_/A _8778_/X _8805_/A vssd1 vssd1 vccd1 vccd1 _8781_/B sky130_fd_sc_hd__o2bb2a_1
X_7800_ _9903_/Q vssd1 vssd1 vccd1 vccd1 _7801_/A sky130_fd_sc_hd__inv_2
X_5992_ _5992_/A vssd1 vssd1 vccd1 vccd1 _5992_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7731_ _7711_/X _7731_/B _7731_/C _7731_/D vssd1 vssd1 vccd1 vccd1 _7773_/B sky130_fd_sc_hd__and4b_1
XFILLER_64_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4943_ _4951_/A vssd1 vssd1 vccd1 vccd1 _4943_/X sky130_fd_sc_hd__buf_1
XFILLER_177_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7662_ _7810_/A _7805_/A vssd1 vssd1 vccd1 vccd1 _7663_/B sky130_fd_sc_hd__or2_1
X_6613_ _6971_/A _7005_/B _6969_/A _7006_/B vssd1 vssd1 vccd1 vccd1 _6613_/X sky130_fd_sc_hd__o22a_1
X_9401_ _9400_/X _7490_/A _9506_/S vssd1 vssd1 vccd1 vccd1 _9401_/X sky130_fd_sc_hd__mux2_1
X_4874_ _9745_/Q _4870_/X _9893_/Q _4871_/X _4873_/X vssd1 vssd1 vccd1 vccd1 _9893_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7593_ _7593_/A _7593_/B vssd1 vssd1 vccd1 vccd1 _7594_/B sky130_fd_sc_hd__or2_1
X_9332_ _9779_/Q _9331_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9332_/X sky130_fd_sc_hd__mux2_1
X_6544_ _6547_/A _6544_/B vssd1 vssd1 vccd1 vccd1 _6544_/Y sky130_fd_sc_hd__nor2_1
X_6475_ _6369_/X _6474_/X _6369_/X _6474_/X vssd1 vssd1 vccd1 vccd1 _6475_/X sky130_fd_sc_hd__o2bb2a_1
X_9263_ _7817_/Y _9758_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9263_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8214_ _8211_/A _8211_/B _6348_/Y _8213_/Y vssd1 vssd1 vccd1 vccd1 _8214_/X sky130_fd_sc_hd__o22a_1
X_5426_ _5426_/A _5426_/B vssd1 vssd1 vccd1 vccd1 _5426_/Y sky130_fd_sc_hd__nor2_1
X_9194_ _6537_/Y _9799_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9548_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8145_ _7819_/A _8117_/X _8144_/X vssd1 vssd1 vccd1 vccd1 _8145_/X sky130_fd_sc_hd__a21o_1
XFILLER_99_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5357_ _5357_/A vssd1 vssd1 vccd1 vccd1 _5358_/B sky130_fd_sc_hd__inv_2
X_8076_ _9548_/Q _8076_/B vssd1 vssd1 vccd1 vccd1 _8077_/B sky130_fd_sc_hd__or2_2
XINSDIODE2_4 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5288_ _5283_/B _5271_/X _5287_/Y _5275_/X _5244_/A vssd1 vssd1 vccd1 vccd1 _5289_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_58_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7027_ _9611_/Q _6691_/B _6756_/A _6610_/Y _7026_/X vssd1 vssd1 vccd1 vccd1 _7027_/X
+ sky130_fd_sc_hd__a41o_2
XFILLER_114_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8978_ _8977_/X _6971_/A _9507_/S vssd1 vssd1 vccd1 vccd1 _8978_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7929_ _7991_/A vssd1 vssd1 vccd1 vccd1 _7956_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_70_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6260_ _9586_/Q _6168_/A _8029_/A _6245_/A vssd1 vssd1 vccd1 vccd1 _6265_/D sky130_fd_sc_hd__a22o_1
XFILLER_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5211_ _5032_/X _5203_/X _9753_/Q _5205_/X _5206_/X vssd1 vssd1 vccd1 vccd1 _9753_/D
+ sky130_fd_sc_hd__a221o_1
X_6191_ _9574_/Q vssd1 vssd1 vccd1 vccd1 _7993_/A sky130_fd_sc_hd__inv_2
X_5142_ _5136_/X _9783_/Q _5138_/X _9210_/X _5140_/X vssd1 vssd1 vccd1 vccd1 _9783_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5073_ _5097_/A vssd1 vssd1 vccd1 vccd1 _5073_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8901_ _8942_/A _8959_/B _8901_/C vssd1 vssd1 vccd1 vccd1 _8901_/X sky130_fd_sc_hd__or3_4
X_9881_ _9895_/CLK _9881_/D vssd1 vssd1 vccd1 vccd1 _9881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8832_ _8832_/A _8904_/A vssd1 vssd1 vccd1 vccd1 _8833_/B sky130_fd_sc_hd__nor2_2
XFILLER_92_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8763_ _8762_/A _8762_/B _8904_/A vssd1 vssd1 vccd1 vccd1 _8763_/X sky130_fd_sc_hd__a21o_1
X_5975_ _5971_/Y _5974_/X _5971_/Y _5974_/X vssd1 vssd1 vccd1 vccd1 _5975_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8694_ _8694_/A vssd1 vssd1 vccd1 vccd1 _8695_/B sky130_fd_sc_hd__inv_2
X_7714_ _9912_/Q vssd1 vssd1 vccd1 vccd1 _7840_/A sky130_fd_sc_hd__inv_2
X_4926_ _9864_/Q _4922_/X _9716_/Q _4920_/X _4923_/X vssd1 vssd1 vccd1 vccd1 _9864_/D
+ sky130_fd_sc_hd__o221a_1
X_7645_ _7652_/B _9707_/Q vssd1 vssd1 vccd1 vccd1 _7645_/Y sky130_fd_sc_hd__nor2b_1
XFILLER_100_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4857_ _5844_/A _7918_/A vssd1 vssd1 vccd1 vccd1 _5976_/A sky130_fd_sc_hd__or2_2
XFILLER_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7576_ _7576_/A _7576_/B vssd1 vssd1 vccd1 vccd1 _7577_/A sky130_fd_sc_hd__or2_1
XFILLER_193_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9315_ _7890_/X _9775_/Q _9327_/S vssd1 vssd1 vccd1 vccd1 _9315_/X sky130_fd_sc_hd__mux2_1
X_4788_ _9921_/Q vssd1 vssd1 vccd1 vccd1 _4788_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6527_ _6529_/A _6527_/B vssd1 vssd1 vccd1 vccd1 _6527_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9246_ _9245_/X _5032_/A _9306_/S vssd1 vssd1 vccd1 vccd1 _9246_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6458_ _6458_/A vssd1 vssd1 vccd1 vccd1 _6458_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6389_ _9771_/Q _8211_/A vssd1 vssd1 vccd1 vccd1 _6390_/B sky130_fd_sc_hd__or2_2
X_9177_ _9176_/X _9783_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9532_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5409_ _5409_/A _5409_/B vssd1 vssd1 vccd1 vccd1 _5409_/Y sky130_fd_sc_hd__nor2_1
X_8128_ _9897_/Q _8128_/B vssd1 vssd1 vccd1 vccd1 _8128_/X sky130_fd_sc_hd__or2_1
XFILLER_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8059_ _4973_/X _8052_/Y _8053_/Y _8058_/Y vssd1 vssd1 vccd1 vccd1 _8059_/X sky130_fd_sc_hd__o22a_1
XFILLER_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5760_ _5757_/Y _5759_/X _5757_/Y _5759_/X vssd1 vssd1 vccd1 vccd1 _9475_/S sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5691_ _6561_/A _5689_/X _9101_/X _5684_/X _5690_/X vssd1 vssd1 vccd1 vccd1 _9674_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_187_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7430_ _7426_/X _7429_/X _7426_/X _7429_/X vssd1 vssd1 vccd1 vccd1 _7430_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _9692_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7361_ _7492_/C _7291_/B _7273_/A _7359_/Y _7360_/X vssd1 vssd1 vccd1 vccd1 _7361_/X
+ sky130_fd_sc_hd__a41o_1
X_6312_ _9799_/Q _9798_/Q _9797_/Q _9796_/Q vssd1 vssd1 vccd1 vccd1 _6315_/B sky130_fd_sc_hd__or4_4
X_9100_ _6020_/X _6022_/X _9896_/Q vssd1 vssd1 vccd1 vccd1 _9100_/X sky130_fd_sc_hd__mux2_1
X_7292_ _7292_/A vssd1 vssd1 vccd1 vccd1 _7292_/Y sky130_fd_sc_hd__inv_2
X_6243_ _6243_/A vssd1 vssd1 vccd1 vccd1 _6265_/A sky130_fd_sc_hd__inv_2
XFILLER_143_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9031_ _7975_/Y _9030_/X _9052_/S vssd1 vssd1 vccd1 vccd1 _9031_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6174_ _9571_/Q vssd1 vssd1 vccd1 vccd1 _7976_/A sky130_fd_sc_hd__inv_2
X_5125_ _4743_/X _9794_/Q _5121_/X _9221_/X _5124_/X vssd1 vssd1 vccd1 vccd1 _9794_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_111_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5056_ _5069_/A _5056_/B vssd1 vssd1 vccd1 vccd1 _9810_/D sky130_fd_sc_hd__nor2_1
XFILLER_65_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9864_ _9874_/CLK _9864_/D vssd1 vssd1 vccd1 vccd1 _9864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8815_ _8765_/A _8786_/X _8788_/B vssd1 vssd1 vccd1 vccd1 _8815_/X sky130_fd_sc_hd__o21a_1
X_9795_ _9929_/CLK _9795_/D vssd1 vssd1 vccd1 vccd1 _9795_/Q sky130_fd_sc_hd__dfxtp_2
X_8746_ _8407_/X _8745_/X _8407_/X _8745_/X vssd1 vssd1 vccd1 vccd1 _8747_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5958_ _5958_/A vssd1 vssd1 vccd1 vccd1 _5958_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_166_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4909_ _9874_/Q _4905_/X _9726_/Q _4903_/X _4906_/X vssd1 vssd1 vccd1 vccd1 _9874_/D
+ sky130_fd_sc_hd__o221a_1
X_8677_ _8677_/A vssd1 vssd1 vccd1 vccd1 _8677_/Y sky130_fd_sc_hd__inv_2
X_5889_ _6713_/A _5884_/X _5032_/A _5885_/X _5875_/X vssd1 vssd1 vccd1 vccd1 _9616_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_138_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7628_ _7070_/A _7070_/B _7071_/B vssd1 vssd1 vccd1 vccd1 _7628_/X sky130_fd_sc_hd__a21bo_1
XFILLER_181_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7559_ _7559_/A _7559_/B vssd1 vssd1 vccd1 vccd1 _7560_/A sky130_fd_sc_hd__and2_1
XFILLER_119_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9229_ _9228_/X _7781_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9229_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6930_ _6923_/Y _6927_/X _6923_/Y _6927_/X vssd1 vssd1 vccd1 vccd1 _6930_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6861_ _6789_/X _6859_/X _6748_/X _6860_/X vssd1 vssd1 vccd1 vccd1 _6861_/X sky130_fd_sc_hd__o211a_1
XFILLER_179_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8600_ _8599_/A _8599_/B _8645_/A vssd1 vssd1 vccd1 vccd1 _8600_/X sky130_fd_sc_hd__a21bo_1
X_9580_ _9833_/CLK _9580_/D vssd1 vssd1 vccd1 vccd1 _9580_/Q sky130_fd_sc_hd__dfxtp_1
X_6792_ _9426_/X vssd1 vssd1 vccd1 vccd1 _6862_/A sky130_fd_sc_hd__clkbuf_2
X_5812_ _6872_/A _5442_/B _5811_/Y _5442_/Y _5811_/A vssd1 vssd1 vccd1 vccd1 _7083_/B
+ sky130_fd_sc_hd__o32a_2
XFILLER_62_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8531_ _8531_/A _8531_/B vssd1 vssd1 vccd1 vccd1 _8531_/Y sky130_fd_sc_hd__nor2_1
X_5743_ _6571_/A _9652_/Q _5442_/Y _5811_/A vssd1 vssd1 vccd1 vccd1 _5744_/A sky130_fd_sc_hd__a22o_1
X_8462_ _8463_/B vssd1 vssd1 vccd1 vccd1 _8462_/Y sky130_fd_sc_hd__inv_2
X_5674_ _5772_/A vssd1 vssd1 vccd1 vccd1 _5674_/X sky130_fd_sc_hd__buf_1
XFILLER_30_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8393_ _9687_/Q vssd1 vssd1 vccd1 vccd1 _8394_/A sky130_fd_sc_hd__inv_2
X_7413_ _7413_/A vssd1 vssd1 vccd1 vccd1 _7415_/A sky130_fd_sc_hd__inv_2
XFILLER_190_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7344_ _7343_/A _7343_/B _7350_/A vssd1 vssd1 vccd1 vccd1 _7347_/A sky130_fd_sc_hd__a21bo_1
XFILLER_190_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7275_ _7160_/A _9471_/X _7156_/A _9472_/X _7274_/Y vssd1 vssd1 vccd1 vccd1 _7276_/B
+ sky130_fd_sc_hd__o41a_1
XFILLER_143_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6226_ _9580_/Q vssd1 vssd1 vccd1 vccd1 _8015_/A sky130_fd_sc_hd__inv_2
X_9014_ _9013_/X _9597_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9014_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6157_ _6155_/X _6156_/Y _6155_/X _6156_/Y vssd1 vssd1 vccd1 vccd1 _6157_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5108_ _9798_/Q vssd1 vssd1 vccd1 vccd1 _5108_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6088_ _6088_/A _6088_/B vssd1 vssd1 vccd1 vccd1 _6088_/X sky130_fd_sc_hd__or2_1
XFILLER_45_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5039_ _5039_/A vssd1 vssd1 vccd1 vccd1 _5039_/X sky130_fd_sc_hd__buf_4
X_9916_ _9916_/CLK _9916_/D vssd1 vssd1 vccd1 vccd1 _9916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9847_ _9907_/CLK _9847_/D vssd1 vssd1 vccd1 vccd1 _9847_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9778_ _9926_/CLK _9778_/D vssd1 vssd1 vccd1 vccd1 _9778_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8729_ _8667_/X _8678_/X _8655_/X _8679_/X vssd1 vssd1 vccd1 vccd1 _8729_/X sky130_fd_sc_hd__o22a_1
XFILLER_15_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput75 _9067_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_163_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput64 _9057_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[19] sky130_fd_sc_hd__clkbuf_2
Xoutput53 _8378_/X vssd1 vssd1 vccd1 vccd1 io_wb_ack_o sky130_fd_sc_hd__clkbuf_2
XFILLER_163_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5390_ _5385_/B _5379_/X _5389_/Y _5327_/A _5364_/A vssd1 vssd1 vccd1 vccd1 _5391_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_99_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7060_ _7060_/A vssd1 vssd1 vccd1 vccd1 _7077_/A sky130_fd_sc_hd__inv_2
X_6011_ _6008_/A _6006_/X _6008_/A _6006_/X vssd1 vssd1 vccd1 vccd1 _6011_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_86_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7962_ _7962_/A _7981_/B vssd1 vssd1 vccd1 vccd1 _7962_/X sky130_fd_sc_hd__or2_1
XFILLER_94_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9701_ _9819_/CLK _9701_/D vssd1 vssd1 vccd1 vccd1 _9701_/Q sky130_fd_sc_hd__dfxtp_1
X_6913_ _6909_/X _6912_/X _6909_/X _6912_/X vssd1 vssd1 vccd1 vccd1 _6913_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7893_ _7897_/B vssd1 vssd1 vccd1 vccd1 _7893_/Y sky130_fd_sc_hd__inv_2
X_9632_ _9750_/CLK _9632_/D vssd1 vssd1 vccd1 vccd1 _9632_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6844_ _9611_/Q _6774_/B _6756_/A _6842_/Y _6843_/X vssd1 vssd1 vccd1 vccd1 _6844_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_35_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9563_ _9761_/CLK _9563_/D vssd1 vssd1 vccd1 vccd1 _9563_/Q sky130_fd_sc_hd__dfxtp_1
X_6775_ _6775_/A vssd1 vssd1 vccd1 vccd1 _6775_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8514_ _8498_/X _8513_/X _8498_/X _8513_/X vssd1 vssd1 vccd1 vccd1 _8514_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_195_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5726_ _9660_/Q vssd1 vssd1 vccd1 vccd1 _5726_/Y sky130_fd_sc_hd__inv_2
X_9494_ _9493_/X _6975_/A _9507_/S vssd1 vssd1 vccd1 vccd1 _9494_/X sky130_fd_sc_hd__mux2_1
X_8445_ _8446_/A vssd1 vssd1 vccd1 vccd1 _8445_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5657_ _9690_/Q _5645_/X _6561_/A _5650_/X _5647_/X vssd1 vssd1 vccd1 vccd1 _9690_/D
+ sky130_fd_sc_hd__o221a_1
X_8376_ _8364_/X _8368_/X _8375_/X _8302_/C vssd1 vssd1 vccd1 vccd1 _8377_/B sky130_fd_sc_hd__o211a_1
X_5588_ _5588_/A _5588_/B vssd1 vssd1 vccd1 vccd1 _5588_/X sky130_fd_sc_hd__and2_1
X_7327_ _7312_/X _7313_/X _7325_/X _7326_/X vssd1 vssd1 vccd1 vccd1 _7327_/X sky130_fd_sc_hd__o22a_1
XFILLER_131_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7258_ _7234_/C _7231_/B _7231_/Y vssd1 vssd1 vccd1 vccd1 _7259_/B sky130_fd_sc_hd__o21ai_1
XFILLER_131_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6209_ _6221_/B _6208_/X _6221_/B _6208_/X vssd1 vssd1 vccd1 vccd1 _6209_/X sky130_fd_sc_hd__a2bb2o_1
X_7189_ _7165_/C _7162_/B _7162_/Y vssd1 vssd1 vccd1 vccd1 _7190_/B sky130_fd_sc_hd__o21ai_1
XFILLER_133_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4890_ _9733_/Q _4865_/X _9881_/Q _4866_/X _4887_/X vssd1 vssd1 vccd1 vccd1 _9881_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6560_ _8389_/B _6558_/B _6559_/Y vssd1 vssd1 vccd1 vccd1 _6560_/X sky130_fd_sc_hd__a21o_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater94 _9294_/S vssd1 vssd1 vccd1 vccd1 _9306_/S sky130_fd_sc_hd__buf_4
X_5511_ _6872_/A vssd1 vssd1 vccd1 vccd1 _6867_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_173_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6491_ _6472_/Y _6480_/A _6478_/Y _6480_/X _6490_/X vssd1 vssd1 vccd1 vccd1 _6491_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8230_ _6331_/A _8229_/X _8227_/Y vssd1 vssd1 vccd1 vccd1 _8230_/X sky130_fd_sc_hd__a21o_1
X_5442_ _5442_/A _5442_/B vssd1 vssd1 vccd1 vccd1 _5442_/Y sky130_fd_sc_hd__nor2_4
XFILLER_172_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8161_ _4802_/A _8105_/Y _8160_/Y vssd1 vssd1 vccd1 vccd1 _8161_/X sky130_fd_sc_hd__o21a_1
X_5373_ _5368_/B _5356_/X _5372_/Y _5331_/A _5364_/X vssd1 vssd1 vccd1 vccd1 _5374_/A
+ sky130_fd_sc_hd__o32a_1
X_8092_ _9558_/Q vssd1 vssd1 vccd1 vccd1 _8092_/Y sky130_fd_sc_hd__inv_2
X_7112_ _9621_/Q vssd1 vssd1 vccd1 vccd1 _7334_/A sky130_fd_sc_hd__inv_2
XFILLER_99_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7043_ _7024_/X _7031_/X _7024_/X _7031_/X vssd1 vssd1 vccd1 vccd1 _7060_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8994_ _8993_/X _6343_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _8994_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7945_ _8606_/A vssd1 vssd1 vccd1 vccd1 _8875_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7876_ _7709_/X _7871_/Y _7679_/B vssd1 vssd1 vccd1 vccd1 _7876_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_82_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9615_ _9656_/CLK _9615_/D vssd1 vssd1 vccd1 vccd1 _9615_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6827_ _6827_/A vssd1 vssd1 vccd1 vccd1 _6829_/A sky130_fd_sc_hd__inv_2
X_9546_ _9916_/CLK _9546_/D vssd1 vssd1 vccd1 vccd1 _9546_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6758_ _6755_/A _9094_/X _6760_/A _9095_/X _6757_/Y vssd1 vssd1 vccd1 vccd1 _6759_/B
+ sky130_fd_sc_hd__o41a_1
XFILLER_148_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9477_ _8560_/Y _8559_/B _9477_/S vssd1 vssd1 vccd1 vccd1 _9477_/X sky130_fd_sc_hd__mux2_2
XFILLER_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6689_ _6676_/X _6686_/X _6687_/X _6688_/X vssd1 vssd1 vccd1 vccd1 _6689_/X sky130_fd_sc_hd__o22a_1
XFILLER_109_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5709_ _5816_/A _5709_/B vssd1 vssd1 vccd1 vccd1 _5710_/A sky130_fd_sc_hd__or2_1
XFILLER_191_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8428_ _8436_/C _8428_/B vssd1 vssd1 vccd1 vccd1 _8440_/A sky130_fd_sc_hd__nand2_1
XFILLER_163_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8359_ _9556_/Q vssd1 vssd1 vccd1 vccd1 _8359_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5991_ _7928_/A _9636_/Q _5704_/C _5981_/Y vssd1 vssd1 vccd1 vccd1 _5992_/A sky130_fd_sc_hd__o22a_1
XFILLER_64_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7730_ _7723_/X _9765_/Q _7726_/X _9757_/Q _7729_/X vssd1 vssd1 vccd1 vccd1 _7731_/D
+ sky130_fd_sc_hd__o221a_1
X_4942_ _9122_/X _4934_/X _9859_/Q _4935_/X _4939_/X vssd1 vssd1 vccd1 vccd1 _9859_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7661_ _9904_/Q _7661_/B vssd1 vssd1 vccd1 vccd1 _7805_/A sky130_fd_sc_hd__or2_1
X_6612_ _7006_/B vssd1 vssd1 vccd1 vccd1 _6612_/Y sky130_fd_sc_hd__inv_2
X_9400_ _9399_/X _8955_/A _9505_/S vssd1 vssd1 vccd1 vccd1 _9400_/X sky130_fd_sc_hd__mux2_1
X_4873_ _5206_/A vssd1 vssd1 vccd1 vccd1 _4873_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7592_ _7592_/A _7592_/B vssd1 vssd1 vccd1 vccd1 _7593_/B sky130_fd_sc_hd__nand2_1
X_9331_ _7908_/X _9779_/Q _9331_/S vssd1 vssd1 vccd1 vccd1 _9331_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6543_ _6547_/A _6543_/B vssd1 vssd1 vccd1 vccd1 _6543_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6474_ _8051_/A _9752_/Q _6359_/Y vssd1 vssd1 vccd1 vccd1 _6474_/X sky130_fd_sc_hd__a21o_1
X_9262_ _9261_/X input47/X _9294_/S vssd1 vssd1 vccd1 vccd1 _9262_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8213_ _8213_/A _8219_/B vssd1 vssd1 vccd1 vccd1 _8213_/Y sky130_fd_sc_hd__nor2_1
XFILLER_133_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5425_ _9355_/X vssd1 vssd1 vccd1 vccd1 _5426_/B sky130_fd_sc_hd__inv_2
XFILLER_160_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9193_ _6535_/Y _9798_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9547_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8144_ _7726_/A _8118_/X _7754_/A _8117_/X _8143_/X vssd1 vssd1 vccd1 vccd1 _8144_/X
+ sky130_fd_sc_hd__o221a_1
X_5356_ _5379_/A vssd1 vssd1 vccd1 vccd1 _5356_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_141_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_5 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8075_ _9547_/Q _8075_/B vssd1 vssd1 vccd1 vccd1 _8076_/B sky130_fd_sc_hd__or2_1
XFILLER_101_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5287_ _9739_/Q _5287_/B vssd1 vssd1 vccd1 vccd1 _5287_/Y sky130_fd_sc_hd__nor2_1
X_7026_ _6978_/A _6971_/B _6683_/A _7005_/B vssd1 vssd1 vccd1 vccd1 _7026_/X sky130_fd_sc_hd__o22a_1
XFILLER_74_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8977_ _8976_/X _7522_/A _9506_/S vssd1 vssd1 vccd1 vccd1 _8977_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7928_ _7928_/A _9503_/S vssd1 vssd1 vccd1 vccd1 _7928_/X sky130_fd_sc_hd__or2_1
XFILLER_70_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7859_ _7861_/A _7854_/Y _7675_/B vssd1 vssd1 vccd1 vccd1 _7859_/Y sky130_fd_sc_hd__o21ai_1
XPHY_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9529_ _9898_/CLK _9529_/D vssd1 vssd1 vccd1 vccd1 _9529_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_149_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5210_ _5029_/X _5203_/X _8236_/A _5205_/X _5206_/X vssd1 vssd1 vccd1 vccd1 _9754_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6190_ _6200_/A _6189_/X _6200_/A _6189_/X vssd1 vssd1 vccd1 vccd1 _6190_/Y sky130_fd_sc_hd__a2bb2oi_1
X_5141_ _5136_/X _9784_/Q _5138_/X _9211_/X _5140_/X vssd1 vssd1 vccd1 vccd1 _9784_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5072_ _9838_/Q vssd1 vssd1 vccd1 vccd1 _5072_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8900_ _8751_/X _8866_/X _8867_/X _8868_/X vssd1 vssd1 vccd1 vccd1 _8900_/X sky130_fd_sc_hd__o22a_1
X_9880_ _9895_/CLK _9880_/D vssd1 vssd1 vccd1 vccd1 _9880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8831_ _8825_/X _8830_/X _8825_/X _8830_/X vssd1 vssd1 vccd1 vccd1 _8903_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_37_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8762_ _8762_/A _8762_/B vssd1 vssd1 vccd1 vccd1 _8904_/A sky130_fd_sc_hd__nor2_2
XFILLER_80_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5974_ _9521_/D _5972_/Y _5973_/Y _9521_/Q vssd1 vssd1 vccd1 vccd1 _5974_/X sky130_fd_sc_hd__a22o_1
X_7713_ _7835_/A vssd1 vssd1 vccd1 vccd1 _7713_/X sky130_fd_sc_hd__buf_2
X_8693_ _8642_/X _8692_/X _8642_/X _8692_/X vssd1 vssd1 vccd1 vccd1 _8694_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4925_ _9865_/Q _4922_/X _9717_/Q _4920_/X _4923_/X vssd1 vssd1 vccd1 vccd1 _9865_/D
+ sky130_fd_sc_hd__o221a_1
X_7644_ _7644_/A vssd1 vssd1 vccd1 vccd1 _7652_/B sky130_fd_sc_hd__buf_1
X_4856_ input5/X input4/X _4856_/C _4856_/D vssd1 vssd1 vccd1 vccd1 _7918_/A sky130_fd_sc_hd__or4_4
XFILLER_60_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7575_ _7201_/A _7384_/B _7487_/C _7101_/X vssd1 vssd1 vccd1 vccd1 _7576_/B sky130_fd_sc_hd__o22a_1
XFILLER_193_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4787_ _9310_/X _4782_/X _4786_/X _4784_/X _4778_/X vssd1 vssd1 vccd1 vccd1 _9922_/D
+ sky130_fd_sc_hd__o221a_1
X_9314_ _9313_/X input34/X _9334_/S vssd1 vssd1 vccd1 vccd1 _9314_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6526_ _6529_/A _6526_/B vssd1 vssd1 vccd1 vccd1 _6526_/Y sky130_fd_sc_hd__nor2_1
XFILLER_180_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9245_ _9244_/X _7799_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9245_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6457_ _6463_/A _6463_/B _6454_/X _6466_/C _6466_/B vssd1 vssd1 vccd1 vccd1 _6458_/A
+ sky130_fd_sc_hd__o311a_1
X_6388_ _9770_/Q _8213_/A vssd1 vssd1 vccd1 vccd1 _8211_/A sky130_fd_sc_hd__or2_2
X_9176_ _9846_/Q _6482_/X _9178_/S vssd1 vssd1 vccd1 vccd1 _9176_/X sky130_fd_sc_hd__mux2_1
X_5408_ _9342_/X vssd1 vssd1 vccd1 vccd1 _5409_/B sky130_fd_sc_hd__inv_2
X_8127_ _8056_/A _9529_/Q _8057_/B vssd1 vssd1 vccd1 vccd1 _8128_/B sky130_fd_sc_hd__a21oi_1
XFILLER_161_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5339_ _5339_/A vssd1 vssd1 vccd1 vccd1 _5692_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8058_ _6365_/Y _9530_/Q _8057_/Y vssd1 vssd1 vccd1 vccd1 _8058_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_125_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7009_ _6986_/X _7008_/X _6986_/X _7008_/X vssd1 vssd1 vccd1 vccd1 _7009_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_71_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5690_ _5772_/A vssd1 vssd1 vccd1 vccd1 _5690_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_187_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7360_ _7195_/A _7222_/B _7156_/A _7359_/A vssd1 vssd1 vccd1 vccd1 _7360_/X sky130_fd_sc_hd__o22a_1
XFILLER_190_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6311_ _9795_/Q _9794_/Q _9793_/Q _9792_/Q vssd1 vssd1 vccd1 vccd1 _6315_/A sky130_fd_sc_hd__or4_4
X_7291_ _9622_/Q _7291_/B _7302_/A vssd1 vssd1 vccd1 vccd1 _7292_/A sky130_fd_sc_hd__and3_1
X_6242_ _8021_/A _6245_/A _9583_/Q _6168_/A vssd1 vssd1 vccd1 vccd1 _6243_/A sky130_fd_sc_hd__o22a_1
XFILLER_115_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9030_ _7976_/Y _9603_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9030_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6173_ _6176_/A _6172_/X _6176_/A _6172_/X vssd1 vssd1 vccd1 vccd1 _6173_/X sky130_fd_sc_hd__a2bb2o_1
X_5124_ _5165_/A vssd1 vssd1 vccd1 vccd1 _5124_/X sky130_fd_sc_hd__buf_1
XFILLER_97_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5055_ _5045_/X _6316_/B _5054_/Y _5050_/X vssd1 vssd1 vccd1 vccd1 _5056_/B sky130_fd_sc_hd__o22a_1
XFILLER_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9863_ _9930_/CLK _9863_/D vssd1 vssd1 vccd1 vccd1 _9863_/Q sky130_fd_sc_hd__dfxtp_1
X_8814_ _8799_/X _8813_/Y _8799_/X _8813_/Y vssd1 vssd1 vccd1 vccd1 _8814_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9794_ _9929_/CLK _9794_/D vssd1 vssd1 vccd1 vccd1 _9794_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8745_ _8384_/A _6578_/A _8384_/Y vssd1 vssd1 vccd1 vccd1 _8745_/X sky130_fd_sc_hd__a21o_1
X_5957_ _9146_/X _5951_/X _9570_/Q _5952_/X vssd1 vssd1 vccd1 vccd1 _9570_/D sky130_fd_sc_hd__a22o_1
X_8676_ _8674_/Y _8715_/B _8674_/Y _8715_/B vssd1 vssd1 vccd1 vccd1 _8677_/A sky130_fd_sc_hd__a2bb2o_1
X_4908_ _9875_/Q _4905_/X _9727_/Q _4903_/X _4906_/X vssd1 vssd1 vccd1 vccd1 _9875_/D
+ sky130_fd_sc_hd__o221a_1
X_5888_ _9616_/Q vssd1 vssd1 vccd1 vccd1 _6713_/A sky130_fd_sc_hd__clkbuf_2
X_7627_ _7594_/A _7594_/B _7595_/B vssd1 vssd1 vccd1 vccd1 _7627_/X sky130_fd_sc_hd__a21bo_1
X_4839_ _9246_/X _4834_/X _8123_/A _4836_/X _4830_/X vssd1 vssd1 vccd1 vccd1 _9902_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_181_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7558_ _7558_/A _7558_/B vssd1 vssd1 vccd1 vccd1 _7559_/B sky130_fd_sc_hd__nand2_1
X_6509_ _9803_/Q _6541_/B _9804_/Q _6543_/B _6508_/X vssd1 vssd1 vccd1 vccd1 _6509_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_107_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7489_ _7197_/A _7488_/A _7204_/X _7200_/A _7500_/A vssd1 vssd1 vccd1 vccd1 _7489_/X
+ sky130_fd_sc_hd__a32o_1
X_9228_ _9749_/Q _9227_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9228_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9159_ _6249_/X input28/X _9170_/S vssd1 vssd1 vccd1 vccd1 _9159_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6860_ _6763_/X _6766_/X _6767_/X _6788_/X vssd1 vssd1 vccd1 vccd1 _6860_/X sky130_fd_sc_hd__o22a_1
X_5811_ _5811_/A vssd1 vssd1 vccd1 vccd1 _5811_/Y sky130_fd_sc_hd__inv_2
X_6791_ _9425_/X vssd1 vssd1 vccd1 vccd1 _6868_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8530_ _8528_/X _8529_/X _8528_/X _8529_/X vssd1 vssd1 vccd1 vccd1 _8530_/X sky130_fd_sc_hd__a2bb2o_1
X_5742_ _9669_/Q _9652_/Q _9669_/Q _9652_/Q vssd1 vssd1 vccd1 vccd1 _5811_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_62_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8461_ _8460_/A _8460_/B _8531_/A vssd1 vssd1 vccd1 vccd1 _8463_/B sky130_fd_sc_hd__a21oi_4
X_5673_ _5790_/A vssd1 vssd1 vccd1 vccd1 _5772_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8392_ _9688_/Q _6564_/X _9688_/Q _6564_/X vssd1 vssd1 vccd1 vccd1 _8392_/X sky130_fd_sc_hd__a2bb2o_1
X_7412_ _7395_/X _7396_/X _7395_/X _7396_/X vssd1 vssd1 vccd1 vccd1 _7413_/A sky130_fd_sc_hd__a2bb2o_1
X_7343_ _7343_/A _7343_/B vssd1 vssd1 vccd1 vccd1 _7350_/A sky130_fd_sc_hd__or2_1
XFILLER_190_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7274_ _7277_/C _7274_/B vssd1 vssd1 vccd1 vccd1 _7274_/Y sky130_fd_sc_hd__nand2_1
X_9013_ _9565_/Q _9896_/Q _9013_/S vssd1 vssd1 vccd1 vccd1 _9013_/X sky130_fd_sc_hd__mux2_1
X_6225_ _6224_/A _6224_/B _6232_/A vssd1 vssd1 vccd1 vccd1 _6225_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_106_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6156_ _7949_/A _6143_/X _6152_/X vssd1 vssd1 vccd1 vccd1 _6156_/Y sky130_fd_sc_hd__o21ai_1
X_5107_ _5115_/A _5107_/B vssd1 vssd1 vccd1 vccd1 _9799_/D sky130_fd_sc_hd__nor2_1
X_6087_ _6087_/A vssd1 vssd1 vccd1 vccd1 _6088_/B sky130_fd_sc_hd__inv_2
X_5038_ _9814_/Q _5028_/X _4860_/X _5030_/X _5036_/X vssd1 vssd1 vccd1 vccd1 _9814_/D
+ sky130_fd_sc_hd__o221a_1
X_9915_ _9915_/CLK _9915_/D vssd1 vssd1 vccd1 vccd1 _9915_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9846_ _9907_/CLK _9846_/D vssd1 vssd1 vccd1 vccd1 _9846_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9777_ _9903_/CLK _9777_/D vssd1 vssd1 vccd1 vccd1 _9777_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_202_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8728_ _8719_/X _8727_/X _8719_/X _8727_/X vssd1 vssd1 vccd1 vccd1 _8728_/X sky130_fd_sc_hd__a2bb2o_1
X_6989_ _6989_/A _6978_/X vssd1 vssd1 vccd1 vccd1 _6989_/X sky130_fd_sc_hd__or2b_1
XFILLER_15_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8659_ _8823_/A _8656_/X _8702_/C _8658_/X vssd1 vssd1 vccd1 vccd1 _8659_/X sky130_fd_sc_hd__a31o_1
XFILLER_178_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput76 _9510_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[2] sky130_fd_sc_hd__clkbuf_2
Xoutput65 _9509_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[1] sky130_fd_sc_hd__clkbuf_2
Xoutput54 _9508_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_163_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _9634_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6010_ _6008_/A _6008_/B _6009_/Y vssd1 vssd1 vccd1 vccd1 _6010_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7961_ _8800_/A vssd1 vssd1 vccd1 vccd1 _8958_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7892_ _7892_/A _7892_/B vssd1 vssd1 vccd1 vccd1 _7897_/B sky130_fd_sc_hd__or2_1
X_9700_ _9819_/CLK _9700_/D vssd1 vssd1 vccd1 vccd1 _9700_/Q sky130_fd_sc_hd__dfxtp_1
X_6912_ _6911_/A _6911_/B _6911_/X vssd1 vssd1 vccd1 vccd1 _6912_/X sky130_fd_sc_hd__a21bo_1
XFILLER_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9631_ _9750_/CLK _9631_/D vssd1 vssd1 vccd1 vccd1 _9631_/Q sky130_fd_sc_hd__dfxtp_1
X_6843_ _6642_/A _6705_/B _6760_/A _6842_/A vssd1 vssd1 vccd1 vccd1 _6843_/X sky130_fd_sc_hd__o22a_1
XFILLER_50_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9562_ _9924_/CLK _9562_/D vssd1 vssd1 vccd1 vccd1 _9562_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6774_ _9614_/Q _6774_/B _6785_/A vssd1 vssd1 vccd1 vccd1 _6775_/A sky130_fd_sc_hd__and3_1
X_8513_ _8479_/A _8479_/B _8512_/A _8479_/Y _8512_/Y vssd1 vssd1 vccd1 vccd1 _8513_/X
+ sky130_fd_sc_hd__o32a_1
X_5725_ _5725_/A vssd1 vssd1 vccd1 vccd1 _8386_/B sky130_fd_sc_hd__clkbuf_2
X_9493_ _9492_/X _7497_/A _9506_/S vssd1 vssd1 vccd1 vccd1 _9493_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8444_ _8399_/X _8446_/B _8399_/X _8446_/B vssd1 vssd1 vccd1 vccd1 _8444_/X sky130_fd_sc_hd__a2bb2o_1
X_5656_ _9674_/Q vssd1 vssd1 vccd1 vccd1 _6561_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_175_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8375_ _8375_/A _8375_/B _8375_/C _8375_/D vssd1 vssd1 vccd1 vccd1 _8375_/X sky130_fd_sc_hd__or4_4
X_5587_ _5587_/A vssd1 vssd1 vccd1 vccd1 _5587_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7326_ _7312_/X _7313_/X _7312_/X _7313_/X vssd1 vssd1 vccd1 vccd1 _7326_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_89_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7257_ _7245_/A _7245_/B _7427_/A vssd1 vssd1 vccd1 vccd1 _7260_/A sky130_fd_sc_hd__a21o_1
XFILLER_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6208_ _9575_/Q _6171_/X _6199_/A _6204_/A vssd1 vssd1 vccd1 vccd1 _6208_/X sky130_fd_sc_hd__a22o_1
X_7188_ _7176_/A _7176_/B _7502_/A vssd1 vssd1 vccd1 vccd1 _7191_/A sky130_fd_sc_hd__a21o_1
XFILLER_58_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6139_ _6139_/A vssd1 vssd1 vccd1 vccd1 _6140_/A sky130_fd_sc_hd__buf_2
XFILLER_58_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9829_ _9916_/CLK _9829_/D vssd1 vssd1 vccd1 vccd1 _9829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater95 _9282_/S vssd1 vssd1 vccd1 vccd1 _9294_/S sky130_fd_sc_hd__buf_4
X_5510_ _5435_/X _5450_/X _5435_/X _5450_/X vssd1 vssd1 vccd1 vccd1 _5510_/X sky130_fd_sc_hd__a2bb2o_4
X_6490_ _6304_/Y _6482_/X _6494_/A _6488_/X _6489_/X vssd1 vssd1 vccd1 vccd1 _6490_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5441_ _9651_/Q vssd1 vssd1 vccd1 vccd1 _5442_/B sky130_fd_sc_hd__inv_2
XFILLER_172_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8160_ _7692_/X _8106_/X _8159_/Y vssd1 vssd1 vccd1 vccd1 _8160_/Y sky130_fd_sc_hd__o21bai_1
X_5372_ _9724_/Q _5372_/B vssd1 vssd1 vccd1 vccd1 _5372_/Y sky130_fd_sc_hd__nor2_1
X_8091_ _8048_/Y _8087_/Y _8089_/X vssd1 vssd1 vccd1 vccd1 _8091_/X sky130_fd_sc_hd__o21a_1
XFILLER_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7111_ _7110_/A _7110_/B _7120_/B vssd1 vssd1 vccd1 vccd1 _7111_/X sky130_fd_sc_hd__a21bo_1
XFILLER_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7042_ _7021_/X _7032_/X _7021_/X _7032_/X vssd1 vssd1 vccd1 vccd1 _7059_/A sky130_fd_sc_hd__a2bb2o_1
X_8993_ _6316_/C _7902_/A _9480_/S vssd1 vssd1 vccd1 vccd1 _8993_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7944_ _9631_/Q vssd1 vssd1 vccd1 vccd1 _8606_/A sky130_fd_sc_hd__inv_2
XFILLER_208_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7875_ _7728_/X _7873_/B _7839_/X _7874_/Y vssd1 vssd1 vccd1 vccd1 _7875_/Y sky130_fd_sc_hd__a211oi_2
XPHY_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9614_ _9656_/CLK _9614_/D vssd1 vssd1 vccd1 vccd1 _9614_/Q sky130_fd_sc_hd__dfxtp_2
X_6826_ _6808_/X _6809_/X _6808_/X _6809_/X vssd1 vssd1 vccd1 vccd1 _6827_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9545_ _9916_/CLK _9545_/D vssd1 vssd1 vccd1 vccd1 _9545_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6757_ _6760_/C _6757_/B vssd1 vssd1 vccd1 vccd1 _6757_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5708_ _5917_/B _5708_/B _5862_/A vssd1 vssd1 vccd1 vccd1 _5709_/B sky130_fd_sc_hd__or3_1
X_9476_ _8646_/X _8644_/A _9490_/S vssd1 vssd1 vccd1 vccd1 _9476_/X sky130_fd_sc_hd__mux2_1
X_6688_ _6676_/X _6686_/X _6676_/X _6686_/X vssd1 vssd1 vccd1 vccd1 _6688_/X sky130_fd_sc_hd__a2bb2o_1
X_8427_ _8427_/A vssd1 vssd1 vccd1 vccd1 _8427_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5639_ _9697_/Q _5631_/X _6593_/A _5635_/X _5632_/X vssd1 vssd1 vccd1 vccd1 _9697_/D
+ sky130_fd_sc_hd__o221a_1
X_8358_ _7709_/X _9553_/Q _8174_/A _9560_/Q vssd1 vssd1 vccd1 vccd1 _8363_/B sky130_fd_sc_hd__a22o_1
XFILLER_191_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7309_ _9474_/X vssd1 vssd1 vccd1 vccd1 _7379_/A sky130_fd_sc_hd__clkbuf_2
X_8289_ _4794_/A _8214_/X _8288_/X vssd1 vssd1 vccd1 vccd1 _8289_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5990_ _5989_/A _5989_/B _5989_/X vssd1 vssd1 vccd1 vccd1 _5990_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4941_ _9123_/X _4934_/X _9860_/Q _4935_/X _4939_/X vssd1 vssd1 vccd1 vccd1 _9860_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_52_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7660_ _9903_/Q _7795_/A vssd1 vssd1 vccd1 vccd1 _7661_/B sky130_fd_sc_hd__or2_1
X_4872_ _5214_/A vssd1 vssd1 vccd1 vccd1 _5206_/A sky130_fd_sc_hd__clkbuf_4
X_6611_ _9462_/X vssd1 vssd1 vccd1 vccd1 _7006_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_60_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9330_ _9329_/X input39/X _9334_/S vssd1 vssd1 vccd1 vccd1 _9330_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7591_ _7591_/A vssd1 vssd1 vccd1 vccd1 _7592_/B sky130_fd_sc_hd__inv_2
X_6542_ _6542_/A vssd1 vssd1 vccd1 vccd1 _6547_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6473_ _9787_/Q _6521_/B vssd1 vssd1 vccd1 vccd1 _6480_/A sky130_fd_sc_hd__nor2_1
X_9261_ _9260_/X _7816_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9261_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8212_ _6390_/B _8211_/B _6413_/Y _8211_/Y vssd1 vssd1 vccd1 vccd1 _8212_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_118_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9192_ _6534_/Y _9797_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9546_/D sky130_fd_sc_hd__mux2_1
X_5424_ _9357_/X vssd1 vssd1 vccd1 vccd1 _5426_/A sky130_fd_sc_hd__inv_2
XFILLER_133_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8143_ _7726_/A _8118_/X _8142_/Y vssd1 vssd1 vccd1 vccd1 _8143_/X sky130_fd_sc_hd__a21o_1
XFILLER_160_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5355_ _5355_/A vssd1 vssd1 vccd1 vccd1 _9728_/D sky130_fd_sc_hd__inv_2
XINSDIODE2_6 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8074_ _9546_/Q _8074_/B vssd1 vssd1 vccd1 vccd1 _8075_/B sky130_fd_sc_hd__or2_1
XFILLER_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5286_ _5286_/A vssd1 vssd1 vccd1 vccd1 _5287_/B sky130_fd_sc_hd__inv_2
XFILLER_87_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7025_ _6938_/X _6957_/Y _6938_/X _6957_/Y vssd1 vssd1 vccd1 vccd1 _7025_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8976_ _8975_/X _8958_/A _9505_/S vssd1 vssd1 vccd1 vccd1 _8976_/X sky130_fd_sc_hd__mux2_1
X_7927_ _8829_/A vssd1 vssd1 vccd1 vccd1 _8935_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_130_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7858_ _7692_/X _7856_/B _7839_/X _7857_/Y vssd1 vssd1 vccd1 vccd1 _7858_/Y sky130_fd_sc_hd__a211oi_2
XPHY_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6809_ _6795_/X _6796_/X _6795_/X _6796_/X vssd1 vssd1 vccd1 vccd1 _6809_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7789_ _7793_/B vssd1 vssd1 vccd1 vccd1 _7789_/Y sky130_fd_sc_hd__inv_2
XPHY_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9528_ _9907_/CLK _9528_/D vssd1 vssd1 vccd1 vccd1 _9528_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9459_ _9803_/Q _9920_/Q _9480_/S vssd1 vssd1 vccd1 vccd1 _9459_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5140_ _5165_/A vssd1 vssd1 vccd1 vccd1 _5140_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5071_ _9806_/Q vssd1 vssd1 vccd1 vccd1 _6317_/B sky130_fd_sc_hd__inv_2
XFILLER_111_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8830_ _8827_/Y _8829_/X _8827_/Y _8829_/X vssd1 vssd1 vccd1 vccd1 _8830_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8761_ _8760_/A _8760_/B _8832_/A vssd1 vssd1 vccd1 vccd1 _8762_/B sky130_fd_sc_hd__a21o_1
X_5973_ _9521_/D vssd1 vssd1 vccd1 vccd1 _5973_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7712_ _9911_/Q vssd1 vssd1 vccd1 vccd1 _7835_/A sky130_fd_sc_hd__inv_2
X_4924_ _9866_/Q _4922_/X _9718_/Q _4920_/X _4923_/X vssd1 vssd1 vccd1 vccd1 _9866_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_40_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8692_ _8683_/X _8691_/X _8683_/X _8691_/X vssd1 vssd1 vccd1 vccd1 _8692_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7643_ _7643_/A _7648_/B vssd1 vssd1 vccd1 vccd1 _7643_/Y sky130_fd_sc_hd__nor2_1
X_4855_ _4855_/A _4855_/B vssd1 vssd1 vccd1 vccd1 _4856_/D sky130_fd_sc_hd__nand2_1
X_4786_ _9922_/Q vssd1 vssd1 vccd1 vccd1 _4786_/X sky130_fd_sc_hd__buf_2
XFILLER_119_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7574_ _7346_/A _7346_/B _7347_/B vssd1 vssd1 vccd1 vccd1 _7592_/A sky130_fd_sc_hd__a21bo_1
X_9313_ _9312_/X _7888_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9313_/X sky130_fd_sc_hd__mux2_1
X_6525_ _6529_/A _6525_/B vssd1 vssd1 vccd1 vccd1 _6525_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9244_ _9753_/Q _9243_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9244_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6456_ _6456_/A _6456_/B vssd1 vssd1 vccd1 vccd1 _6466_/B sky130_fd_sc_hd__or2_2
X_9175_ _9174_/X _9782_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9531_/D sky130_fd_sc_hd__mux2_1
X_6387_ _9769_/Q _6418_/A vssd1 vssd1 vccd1 vccd1 _8213_/A sky130_fd_sc_hd__or2_4
X_5407_ _9344_/X vssd1 vssd1 vccd1 vccd1 _5409_/A sky130_fd_sc_hd__inv_2
X_8126_ _8059_/X _8125_/X _8059_/X _8125_/X vssd1 vssd1 vccd1 vccd1 _8126_/Y sky130_fd_sc_hd__o2bb2ai_1
X_5338_ _9731_/Q vssd1 vssd1 vccd1 vccd1 _5338_/Y sky130_fd_sc_hd__inv_2
X_8057_ _8057_/A _8057_/B vssd1 vssd1 vccd1 vccd1 _8057_/Y sky130_fd_sc_hd__nor2_2
XFILLER_114_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7008_ _7004_/Y _7007_/X _7004_/Y _7007_/X vssd1 vssd1 vccd1 vccd1 _7008_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5269_ _5264_/B _5224_/X _5268_/Y _4853_/X _5248_/A vssd1 vssd1 vccd1 vccd1 _5270_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_87_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8959_ _8959_/A _8959_/B vssd1 vssd1 vccd1 vccd1 _8959_/Y sky130_fd_sc_hd__nor2_1
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6310_ _4960_/X _6309_/Y _4973_/X _6304_/Y vssd1 vssd1 vccd1 vccd1 _6310_/X sky130_fd_sc_hd__a22o_1
XFILLER_128_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7290_ _7290_/A _7359_/A vssd1 vssd1 vccd1 vccd1 _7302_/A sky130_fd_sc_hd__or2_1
X_6241_ _6241_/A vssd1 vssd1 vccd1 vccd1 _6245_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6172_ _9569_/Q _6171_/X _6159_/X _6161_/Y vssd1 vssd1 vccd1 vccd1 _6172_/X sky130_fd_sc_hd__a22o_1
X_5123_ _5790_/A vssd1 vssd1 vccd1 vccd1 _5165_/A sky130_fd_sc_hd__buf_2
X_5054_ _9842_/Q vssd1 vssd1 vccd1 vccd1 _5054_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9862_ _9895_/CLK _9862_/D vssd1 vssd1 vccd1 vccd1 _9862_/Q sky130_fd_sc_hd__dfxtp_2
X_8813_ _8812_/A _8812_/B _8812_/Y vssd1 vssd1 vccd1 vccd1 _8813_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_25_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9793_ _9929_/CLK _9793_/D vssd1 vssd1 vccd1 vccd1 _9793_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8744_ _8743_/A _8743_/B _8793_/A vssd1 vssd1 vccd1 vccd1 _8744_/X sky130_fd_sc_hd__a21bo_1
XFILLER_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5956_ _9147_/X _5951_/X _9571_/Q _5952_/X vssd1 vssd1 vccd1 vccd1 _9571_/D sky130_fd_sc_hd__a22o_1
X_8675_ _8766_/C _8626_/X _8627_/X _8631_/X vssd1 vssd1 vccd1 vccd1 _8715_/B sky130_fd_sc_hd__o22ai_2
X_5887_ _9617_/Q _5884_/X _5029_/A _5885_/X _5875_/X vssd1 vssd1 vccd1 vccd1 _9617_/D
+ sky130_fd_sc_hd__o221a_1
X_4907_ _9876_/Q _4905_/X _9728_/Q _4903_/X _4906_/X vssd1 vssd1 vccd1 vccd1 _9876_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_166_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4838_ _9902_/Q vssd1 vssd1 vccd1 vccd1 _8123_/A sky130_fd_sc_hd__clkbuf_2
X_7626_ _7071_/A _7071_/B _7072_/B vssd1 vssd1 vccd1 vccd1 _7626_/X sky130_fd_sc_hd__a21bo_1
XFILLER_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4769_ _9927_/Q vssd1 vssd1 vccd1 vccd1 _7684_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7557_ _7558_/A _7558_/B vssd1 vssd1 vccd1 vccd1 _7559_/A sky130_fd_sc_hd__or2_1
XFILLER_181_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6508_ _9802_/Q _6540_/B _9803_/Q _6541_/B _6507_/X vssd1 vssd1 vccd1 vccd1 _6508_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7488_ _7488_/A vssd1 vssd1 vccd1 vccd1 _7500_/A sky130_fd_sc_hd__inv_2
X_9227_ _7781_/B _9749_/Q _9327_/S vssd1 vssd1 vccd1 vccd1 _9227_/X sky130_fd_sc_hd__mux2_1
X_6439_ _6335_/A _8231_/A _6435_/Y vssd1 vssd1 vccd1 vccd1 _6528_/B sky130_fd_sc_hd__a21oi_4
X_9158_ _6239_/X input26/X _9170_/S vssd1 vssd1 vccd1 vccd1 _9158_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8109_ _9545_/Q _8073_/B _8074_/B vssd1 vssd1 vccd1 vccd1 _8109_/X sky130_fd_sc_hd__a21bo_1
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9089_ _9767_/Q _9088_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9089_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5810_ _9653_/Q _5793_/X _4900_/X _7084_/A _5809_/X vssd1 vssd1 vccd1 vccd1 _9653_/D
+ sky130_fd_sc_hd__o221a_1
X_6790_ _6786_/A _6786_/B _6855_/B vssd1 vssd1 vccd1 vccd1 _6790_/X sky130_fd_sc_hd__a21o_1
X_5741_ _9670_/Q _9653_/Q vssd1 vssd1 vccd1 vccd1 _5741_/Y sky130_fd_sc_hd__nor2_1
X_8460_ _8460_/A _8460_/B vssd1 vssd1 vccd1 vccd1 _8531_/A sky130_fd_sc_hd__nor2_4
XFILLER_148_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5672_ _9668_/Q vssd1 vssd1 vccd1 vccd1 _6804_/C sky130_fd_sc_hd__buf_2
XFILLER_30_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7411_ _7406_/X _7410_/X _7406_/X _7410_/X vssd1 vssd1 vccd1 vccd1 _7443_/A sky130_fd_sc_hd__a2bb2o_1
X_8391_ _9689_/Q _8391_/B vssd1 vssd1 vccd1 vccd1 _8391_/Y sky130_fd_sc_hd__nor2_1
XFILLER_163_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7342_ _7323_/A _7323_/B _7323_/X vssd1 vssd1 vccd1 vccd1 _7343_/B sky130_fd_sc_hd__a21bo_1
X_7273_ _7273_/A _7273_/B _7367_/A vssd1 vssd1 vccd1 vccd1 _7274_/B sky130_fd_sc_hd__and3_1
X_9012_ _9011_/X _9750_/Q _9481_/S vssd1 vssd1 vccd1 vccd1 _9012_/X sky130_fd_sc_hd__mux2_2
XFILLER_89_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6224_ _6224_/A _6224_/B vssd1 vssd1 vccd1 vccd1 _6232_/A sky130_fd_sc_hd__or2_2
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6155_ _9568_/Q _6165_/A _7957_/A _6135_/A vssd1 vssd1 vccd1 vccd1 _6155_/X sky130_fd_sc_hd__a22o_1
X_5106_ _5084_/X _5104_/Y _5105_/Y _5097_/X vssd1 vssd1 vccd1 vccd1 _5107_/B sky130_fd_sc_hd__o22a_1
XFILLER_97_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6086_ _6057_/Y _6066_/A _6076_/A _6049_/Y _6085_/X vssd1 vssd1 vccd1 vccd1 _6087_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_85_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5037_ _9815_/Q _5028_/X _5035_/X _5030_/X _5036_/X vssd1 vssd1 vccd1 vccd1 _9815_/D
+ sky130_fd_sc_hd__o221a_1
X_9914_ _9915_/CLK _9914_/D vssd1 vssd1 vccd1 vccd1 _9914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9845_ _9907_/CLK _9845_/D vssd1 vssd1 vccd1 vccd1 _9845_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9776_ _9898_/CLK _9776_/D vssd1 vssd1 vccd1 vccd1 _9776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8727_ _8810_/A _8727_/B vssd1 vssd1 vccd1 vccd1 _8727_/X sky130_fd_sc_hd__or2_1
X_6988_ _6978_/A _9465_/X _6978_/C _6981_/B vssd1 vssd1 vccd1 vccd1 _6989_/A sky130_fd_sc_hd__o22a_1
XFILLER_25_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5939_ _9160_/X _5937_/X _9584_/Q _5938_/X vssd1 vssd1 vccd1 vccd1 _9584_/D sky130_fd_sc_hd__a22o_1
XFILLER_15_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8658_ _8821_/A _8768_/A _8576_/A _8800_/B vssd1 vssd1 vccd1 vccd1 _8658_/X sky130_fd_sc_hd__o22a_1
XFILLER_166_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8589_ _8589_/A _8589_/B vssd1 vssd1 vccd1 vccd1 _8633_/A sky130_fd_sc_hd__nor2_2
XFILLER_166_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7609_ _7603_/A _7603_/B _7604_/B vssd1 vssd1 vccd1 vccd1 _7609_/X sky130_fd_sc_hd__a21bo_1
XFILLER_147_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput66 _9058_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[20] sky130_fd_sc_hd__clkbuf_2
Xoutput55 _9038_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[10] sky130_fd_sc_hd__clkbuf_2
Xoutput77 _9068_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_88_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_1_clock clkbuf_1_0_1_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7960_ _8773_/A vssd1 vssd1 vccd1 vccd1 _8800_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7891_ _7891_/A vssd1 vssd1 vccd1 vccd1 _7892_/A sky130_fd_sc_hd__clkbuf_2
X_6911_ _6911_/A _6911_/B vssd1 vssd1 vccd1 vccd1 _6911_/X sky130_fd_sc_hd__or2_1
XFILLER_47_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9630_ _9634_/CLK _9630_/D vssd1 vssd1 vccd1 vccd1 _9630_/Q sky130_fd_sc_hd__dfxtp_1
X_6842_ _6842_/A vssd1 vssd1 vccd1 vccd1 _6842_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9561_ _9928_/CLK _9561_/D vssd1 vssd1 vccd1 vccd1 _9561_/Q sky130_fd_sc_hd__dfxtp_1
X_6773_ _6812_/A _6842_/A vssd1 vssd1 vccd1 vccd1 _6785_/A sky130_fd_sc_hd__or2_1
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8512_ _8512_/A vssd1 vssd1 vccd1 vccd1 _8512_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5724_ _9677_/Q vssd1 vssd1 vccd1 vccd1 _5725_/A sky130_fd_sc_hd__inv_2
X_9492_ _9491_/X _8938_/A _9505_/S vssd1 vssd1 vccd1 vccd1 _9492_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5655_ _9691_/Q _5645_/X _8389_/B _5650_/X _5647_/X vssd1 vssd1 vccd1 vccd1 _9691_/D
+ sky130_fd_sc_hd__o221a_1
X_8443_ _8394_/A _8394_/B _8394_/Y vssd1 vssd1 vccd1 vccd1 _8446_/B sky130_fd_sc_hd__a21o_1
XFILLER_191_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8374_ _8374_/A _8374_/B vssd1 vssd1 vccd1 vccd1 _8375_/A sky130_fd_sc_hd__nand2_1
XFILLER_190_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5586_ _5586_/A vssd1 vssd1 vccd1 vccd1 _5586_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7325_ _7314_/X _7315_/X _7323_/X _7324_/X vssd1 vssd1 vccd1 vccd1 _7325_/X sky130_fd_sc_hd__o22a_1
XFILLER_144_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7256_ _7256_/A vssd1 vssd1 vccd1 vccd1 _7427_/A sky130_fd_sc_hd__inv_2
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6207_ _9576_/Q _6167_/A _8001_/A _6201_/A vssd1 vssd1 vccd1 vccd1 _6221_/B sky130_fd_sc_hd__a22o_1
X_7187_ _7187_/A vssd1 vssd1 vccd1 vccd1 _7502_/A sky130_fd_sc_hd__inv_2
XFILLER_131_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6138_ _6241_/A vssd1 vssd1 vccd1 vccd1 _6139_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6069_ _6066_/Y _6068_/A _6066_/A _6068_/Y vssd1 vssd1 vccd1 vccd1 _6069_/X sky130_fd_sc_hd__o22a_1
XFILLER_26_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9828_ _9828_/CLK _9828_/D vssd1 vssd1 vccd1 vccd1 _9828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9759_ _9909_/CLK _9759_/D vssd1 vssd1 vccd1 vccd1 _9759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5440_ _5442_/A vssd1 vssd1 vccd1 vccd1 _6796_/C sky130_fd_sc_hd__buf_2
XFILLER_8_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5371_ _5371_/A vssd1 vssd1 vccd1 vccd1 _5372_/B sky130_fd_sc_hd__inv_2
X_8090_ _8048_/Y _8087_/Y _8088_/Y _9560_/Q _8089_/X vssd1 vssd1 vccd1 vccd1 _8174_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_126_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7110_ _7110_/A _7110_/B vssd1 vssd1 vccd1 vccd1 _7120_/B sky130_fd_sc_hd__or2_1
XFILLER_113_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7041_ _7018_/X _7033_/X _7018_/X _7033_/X vssd1 vssd1 vccd1 vccd1 _7058_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8992_ _8991_/X _9759_/Q _9481_/S vssd1 vssd1 vccd1 vccd1 _8992_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7943_ _7943_/A _9013_/S vssd1 vssd1 vccd1 vccd1 _7943_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7874_ _7877_/B vssd1 vssd1 vccd1 vccd1 _7874_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9613_ _9656_/CLK _9613_/D vssd1 vssd1 vccd1 vccd1 _9613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6825_ _6820_/X _6824_/X _6820_/X _6824_/X vssd1 vssd1 vccd1 vccd1 _6847_/A sky130_fd_sc_hd__a2bb2o_1
X_9544_ _9916_/CLK _9544_/D vssd1 vssd1 vccd1 vccd1 _9544_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6756_ _6756_/A _6756_/B _6851_/A vssd1 vssd1 vccd1 vccd1 _6757_/B sky130_fd_sc_hd__and3_1
XFILLER_10_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5707_ _5707_/A _5707_/B _5707_/C input9/X vssd1 vssd1 vccd1 vccd1 _5708_/B sky130_fd_sc_hd__or4b_4
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6687_ _6622_/A _6622_/B _6622_/Y vssd1 vssd1 vccd1 vccd1 _6687_/X sky130_fd_sc_hd__a21o_1
X_9475_ _7102_/Y _6115_/Y _9475_/S vssd1 vssd1 vccd1 vccd1 _9475_/X sky130_fd_sc_hd__mux2_2
Xclkbuf_leaf_17_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _9519_/CLK sky130_fd_sc_hd__clkbuf_16
X_8426_ _8426_/A _8428_/B vssd1 vssd1 vccd1 vccd1 _8427_/A sky130_fd_sc_hd__or2_1
XFILLER_163_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5638_ _8381_/B vssd1 vssd1 vccd1 vccd1 _6593_/A sky130_fd_sc_hd__clkbuf_2
X_8357_ _8357_/A _8357_/B _8357_/C _8356_/X vssd1 vssd1 vccd1 vccd1 _8363_/A sky130_fd_sc_hd__or4b_4
XFILLER_191_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5569_ _5579_/A _5569_/B vssd1 vssd1 vccd1 vccd1 _9712_/D sky130_fd_sc_hd__nor2_1
XFILLER_151_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7308_ _9473_/X vssd1 vssd1 vccd1 vccd1 _7385_/B sky130_fd_sc_hd__clkbuf_2
X_8288_ _4798_/A _8217_/X _4794_/A _8214_/X _8287_/X vssd1 vssd1 vccd1 vccd1 _8288_/X
+ sky130_fd_sc_hd__a221o_1
X_7239_ _7239_/A vssd1 vssd1 vccd1 vccd1 _7240_/C sky130_fd_sc_hd__inv_2
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4940_ _9124_/X _4934_/X _9861_/Q _4935_/X _4939_/X vssd1 vssd1 vccd1 vccd1 _9861_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_205_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4871_ _4880_/A vssd1 vssd1 vccd1 vccd1 _4871_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6610_ _7005_/B vssd1 vssd1 vccd1 vccd1 _6610_/Y sky130_fd_sc_hd__inv_2
X_7590_ _7201_/A _7101_/X _7576_/B vssd1 vssd1 vccd1 vccd1 _7591_/A sky130_fd_sc_hd__o21ai_1
XFILLER_177_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6541_ _6541_/A _6541_/B vssd1 vssd1 vccd1 vccd1 _6541_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6472_ _6480_/C vssd1 vssd1 vccd1 vccd1 _6472_/Y sky130_fd_sc_hd__inv_2
X_9260_ _9757_/Q _9259_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9260_/X sky130_fd_sc_hd__mux2_1
X_8211_ _8211_/A _8211_/B vssd1 vssd1 vccd1 vccd1 _8211_/Y sky130_fd_sc_hd__nor2_1
XFILLER_145_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9191_ _6533_/Y _9796_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9545_/D sky130_fd_sc_hd__mux2_1
XFILLER_106_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5423_ _5423_/A _5423_/B vssd1 vssd1 vccd1 vccd1 _5423_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8142_ _7769_/A _8119_/Y _8141_/X vssd1 vssd1 vccd1 vccd1 _8142_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5354_ _5347_/B _5313_/X _5353_/Y _5335_/A _5349_/X vssd1 vssd1 vccd1 vccd1 _5355_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_141_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_7 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8073_ _9545_/Q _8073_/B vssd1 vssd1 vccd1 vccd1 _8074_/B sky130_fd_sc_hd__or2_1
X_5285_ _5285_/A vssd1 vssd1 vccd1 vccd1 _9740_/D sky130_fd_sc_hd__inv_2
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7024_ _7022_/X _7023_/X _7022_/X _7023_/X vssd1 vssd1 vccd1 vccd1 _7024_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8975_ _7962_/X _6023_/Y _9504_/S vssd1 vssd1 vccd1 vccd1 _8975_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7926_ _8735_/A vssd1 vssd1 vccd1 vccd1 _8829_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7857_ _7861_/B vssd1 vssd1 vccd1 vccd1 _7857_/Y sky130_fd_sc_hd__inv_2
XPHY_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6808_ _6797_/X _6798_/X _6806_/X _6807_/X vssd1 vssd1 vccd1 vccd1 _6808_/X sky130_fd_sc_hd__o22a_1
XPHY_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7788_ _7788_/A _7788_/B vssd1 vssd1 vccd1 vccd1 _7793_/B sky130_fd_sc_hd__or2_1
XPHY_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9527_ _9861_/CLK _9527_/D vssd1 vssd1 vccd1 vccd1 _9527_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6739_ _6739_/A vssd1 vssd1 vccd1 vccd1 _6910_/A sky130_fd_sc_hd__inv_2
XFILLER_23_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9458_ _7111_/X _5776_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9458_/X sky130_fd_sc_hd__mux2_2
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8409_ _9696_/Q _6596_/Y _8382_/X _8408_/X vssd1 vssd1 vccd1 vccd1 _8409_/X sky130_fd_sc_hd__o22a_1
XFILLER_191_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9389_ _9388_/X _8204_/A _9481_/S vssd1 vssd1 vccd1 vccd1 _9389_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5070_ _5070_/A vssd1 vssd1 vccd1 vccd1 _5092_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8760_ _8760_/A _8760_/B vssd1 vssd1 vccd1 vccd1 _8832_/A sky130_fd_sc_hd__nor2_2
X_5972_ _9521_/Q vssd1 vssd1 vccd1 vccd1 _5972_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7711_ _4832_/X _6469_/Y _7807_/A _9755_/Q _7710_/X vssd1 vssd1 vccd1 vccd1 _7711_/X
+ sky130_fd_sc_hd__a221o_1
X_4923_ _4923_/A vssd1 vssd1 vccd1 vccd1 _4923_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8691_ _5858_/X _8823_/B _8735_/C _8690_/X vssd1 vssd1 vccd1 vccd1 _8691_/X sky130_fd_sc_hd__a31o_1
XFILLER_138_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7642_ _7642_/A _7648_/B vssd1 vssd1 vccd1 vccd1 _7642_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4854_ _5918_/A vssd1 vssd1 vccd1 vccd1 _5816_/A sky130_fd_sc_hd__buf_2
X_4785_ _9314_/X _4782_/X _7680_/A _4784_/X _4778_/X vssd1 vssd1 vccd1 vccd1 _9923_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7573_ _7347_/A _7347_/B _7348_/B vssd1 vssd1 vccd1 vccd1 _7589_/A sky130_fd_sc_hd__a21bo_1
X_9312_ _9774_/Q _9311_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9312_/X sky130_fd_sc_hd__mux2_1
X_6524_ _6550_/A vssd1 vssd1 vccd1 vccd1 _6529_/A sky130_fd_sc_hd__clkbuf_2
X_9243_ _7796_/X _9753_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9243_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6455_ _9792_/Q _6528_/B vssd1 vssd1 vccd1 vccd1 _6466_/C sky130_fd_sc_hd__nand2_2
X_9174_ _9845_/Q _6487_/B _9178_/S vssd1 vssd1 vccd1 vccd1 _9174_/X sky130_fd_sc_hd__mux2_1
X_6386_ _9768_/Q _8215_/A vssd1 vssd1 vccd1 vccd1 _6418_/A sky130_fd_sc_hd__or2_1
X_5406_ _9340_/X _9339_/X _9340_/X _9339_/X vssd1 vssd1 vccd1 vccd1 _5406_/X sky130_fd_sc_hd__a2bb2o_1
X_8125_ _8051_/A _9532_/Q _8051_/Y vssd1 vssd1 vccd1 vccd1 _8125_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5337_ _5337_/A _5344_/A vssd1 vssd1 vccd1 vccd1 _5340_/C sky130_fd_sc_hd__or2_1
X_8056_ _8056_/A _9529_/Q vssd1 vssd1 vccd1 vccd1 _8057_/B sky130_fd_sc_hd__nor2_2
X_5268_ _9743_/Q _5268_/B vssd1 vssd1 vccd1 vccd1 _5268_/Y sky130_fd_sc_hd__nor2_1
X_7007_ _7005_/X _7006_/Y _7005_/X _7006_/Y vssd1 vssd1 vccd1 vccd1 _7007_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_87_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5199_ input18/X _5192_/X _5198_/X _5193_/X _5194_/X vssd1 vssd1 vccd1 vccd1 _9759_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8958_ _8958_/A _8958_/B vssd1 vssd1 vccd1 vccd1 _8958_/X sky130_fd_sc_hd__or2_1
XFILLER_71_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7909_ _7909_/A vssd1 vssd1 vccd1 vccd1 _7909_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8889_ _8379_/X _8410_/X _8379_/X _8410_/X vssd1 vssd1 vccd1 vccd1 _8890_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_70_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6240_ _9583_/Q vssd1 vssd1 vccd1 vccd1 _8021_/A sky130_fd_sc_hd__inv_2
XFILLER_6_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6171_ _6171_/A vssd1 vssd1 vccd1 vccd1 _6171_/X sky130_fd_sc_hd__buf_4
XFILLER_170_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5122_ _4743_/X _9795_/Q _5121_/X _9222_/X _5036_/X vssd1 vssd1 vccd1 vccd1 _9795_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_97_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5053_ _9810_/Q vssd1 vssd1 vccd1 vccd1 _6316_/B sky130_fd_sc_hd__inv_2
XFILLER_97_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9930_ _9930_/CLK _9930_/D vssd1 vssd1 vccd1 vccd1 _9930_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9861_ _9861_/CLK _9861_/D vssd1 vssd1 vccd1 vccd1 _9861_/Q sky130_fd_sc_hd__dfxtp_1
X_8812_ _8812_/A _8812_/B vssd1 vssd1 vccd1 vccd1 _8812_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9792_ _9929_/CLK _9792_/D vssd1 vssd1 vccd1 vccd1 _9792_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8743_ _8743_/A _8743_/B vssd1 vssd1 vccd1 vccd1 _8793_/A sky130_fd_sc_hd__or2_1
XFILLER_80_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5955_ _9148_/X _5951_/X _9572_/Q _5952_/X vssd1 vssd1 vccd1 vccd1 _9572_/D sky130_fd_sc_hd__a22o_1
X_8674_ _8672_/X _8673_/X _8672_/X _8673_/X vssd1 vssd1 vccd1 vccd1 _8674_/Y sky130_fd_sc_hd__a2bb2oi_2
X_5886_ _9618_/Q _5884_/X _5026_/A _5885_/X _5875_/X vssd1 vssd1 vccd1 vccd1 _9618_/D
+ sky130_fd_sc_hd__o221a_1
X_4906_ _4923_/A vssd1 vssd1 vccd1 vccd1 _4906_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4837_ _9250_/X _4834_/X _4835_/X _4836_/X _4830_/X vssd1 vssd1 vccd1 vccd1 _9903_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_138_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7625_ _7595_/A _7595_/B _7596_/B vssd1 vssd1 vccd1 vccd1 _7625_/X sky130_fd_sc_hd__a21bo_1
XFILLER_119_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4768_ _9334_/X _4763_/X _8301_/A _4767_/X _5916_/A vssd1 vssd1 vccd1 vccd1 _9928_/D
+ sky130_fd_sc_hd__o221a_1
X_7556_ _7526_/X _7555_/Y _7526_/X _7555_/Y vssd1 vssd1 vccd1 vccd1 _7558_/B sky130_fd_sc_hd__a2bb2o_1
X_6507_ _9802_/Q _6540_/B _9801_/Q _6539_/B _6506_/Y vssd1 vssd1 vccd1 vccd1 _6507_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_134_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7487_ _7487_/A _9432_/X _7487_/C _7491_/B vssd1 vssd1 vccd1 vccd1 _7488_/A sky130_fd_sc_hd__or4_4
X_9226_ _9225_/X _5041_/A _9334_/S vssd1 vssd1 vccd1 vccd1 _9226_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6438_ _9793_/Q _6529_/B vssd1 vssd1 vccd1 vccd1 _6465_/B sky130_fd_sc_hd__or2_1
XFILLER_161_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9157_ _6235_/Y input25/X _9170_/S vssd1 vssd1 vccd1 vccd1 _9157_/X sky130_fd_sc_hd__mux2_1
X_6369_ _4973_/X _6360_/Y _6363_/Y _6368_/X vssd1 vssd1 vccd1 vccd1 _6369_/X sky130_fd_sc_hd__o22a_1
X_8108_ _9546_/Q _8074_/B _8075_/B vssd1 vssd1 vccd1 vccd1 _8108_/X sky130_fd_sc_hd__a21bo_1
XFILLER_96_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9088_ _7855_/X _9767_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9088_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8039_ _9438_/X _8047_/B vssd1 vssd1 vccd1 vccd1 _8039_/X sky130_fd_sc_hd__and2_1
XFILLER_29_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5740_ _9671_/Q _9654_/Q vssd1 vssd1 vccd1 vccd1 _5740_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_3_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clock/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5671_ _5689_/A vssd1 vssd1 vccd1 vccd1 _5671_/X sky130_fd_sc_hd__buf_1
X_7410_ _7400_/C _7409_/A _7399_/A _7409_/Y vssd1 vssd1 vccd1 vccd1 _7410_/X sky130_fd_sc_hd__a22o_1
XFILLER_163_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8390_ _9690_/Q _6561_/Y _9690_/Q _6561_/Y vssd1 vssd1 vccd1 vccd1 _8390_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_128_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7341_ _7341_/A _7313_/X vssd1 vssd1 vccd1 vccd1 _7343_/A sky130_fd_sc_hd__or2b_1
XFILLER_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7272_ _7317_/A _9472_/X vssd1 vssd1 vccd1 vccd1 _7367_/A sky130_fd_sc_hd__or2_1
X_9011_ _9782_/Q _9899_/Q _9480_/S vssd1 vssd1 vccd1 vccd1 _9011_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6223_ _6203_/A _6221_/X _6203_/B _6222_/X vssd1 vssd1 vccd1 vccd1 _6224_/B sky130_fd_sc_hd__o211a_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6154_ _9568_/Q vssd1 vssd1 vccd1 vccd1 _7957_/A sky130_fd_sc_hd__inv_2
X_5105_ _9831_/Q vssd1 vssd1 vccd1 vccd1 _5105_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6085_ _7990_/A _9646_/Q _6074_/Y _6079_/X vssd1 vssd1 vccd1 vccd1 _6085_/X sky130_fd_sc_hd__o22a_2
X_5036_ _5036_/A vssd1 vssd1 vccd1 vccd1 _5036_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9913_ _9915_/CLK _9913_/D vssd1 vssd1 vccd1 vccd1 _9913_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_38_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9844_ _9907_/CLK _9844_/D vssd1 vssd1 vccd1 vccd1 _9844_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_72_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9775_ _9926_/CLK _9775_/D vssd1 vssd1 vccd1 vccd1 _9775_/Q sky130_fd_sc_hd__dfxtp_1
X_6987_ _6687_/X _6688_/X _6687_/X _6688_/X vssd1 vssd1 vccd1 vccd1 _6987_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8726_ _8958_/A _8725_/B _8725_/C vssd1 vssd1 vccd1 vccd1 _8727_/B sky130_fd_sc_hd__o21a_1
X_5938_ _5938_/A vssd1 vssd1 vccd1 vccd1 _5938_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8657_ _9457_/X vssd1 vssd1 vccd1 vccd1 _8800_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_178_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5869_ _9625_/Q _5865_/X _5029_/X _5866_/X _5867_/X vssd1 vssd1 vccd1 vccd1 _9625_/D
+ sky130_fd_sc_hd__o221a_1
X_8588_ _8586_/X _8628_/A _8586_/X _8628_/A vssd1 vssd1 vccd1 vccd1 _8589_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_166_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7608_ _7080_/A _7080_/B _7081_/B vssd1 vssd1 vccd1 vccd1 _7608_/X sky130_fd_sc_hd__a21bo_1
XFILLER_193_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7539_ _7536_/X _7538_/X _7536_/X _7538_/X vssd1 vssd1 vccd1 vccd1 _7539_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9209_ _9814_/Q _7638_/Y _9528_/Q vssd1 vssd1 vccd1 vccd1 _9209_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput67 _9059_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_134_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput56 _9041_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[11] sky130_fd_sc_hd__clkbuf_2
Xoutput78 _9069_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_88_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7890_ _4780_/X _7681_/B _7889_/Y vssd1 vssd1 vccd1 vccd1 _7890_/X sky130_fd_sc_hd__a21o_1
X_6910_ _6910_/A _6910_/B vssd1 vssd1 vccd1 vccd1 _6911_/B sky130_fd_sc_hd__nor2_1
XFILLER_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6841_ _6839_/X _6840_/X _6839_/X _6840_/X vssd1 vssd1 vccd1 vccd1 _6841_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9560_ _9926_/CLK _9560_/D vssd1 vssd1 vccd1 vccd1 _9560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8511_ _8510_/A _8531_/B _8510_/Y vssd1 vssd1 vccd1 vccd1 _8512_/A sky130_fd_sc_hd__a21oi_2
XFILLER_195_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6772_ _6759_/X _6760_/X _6759_/X _6760_/X vssd1 vssd1 vccd1 vccd1 _6772_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_50_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5723_ _6577_/A _9661_/Q _5721_/A _5722_/Y vssd1 vssd1 vccd1 vccd1 _5723_/X sky130_fd_sc_hd__a22o_1
X_9491_ _7935_/X _5985_/Y _9504_/S vssd1 vssd1 vccd1 vccd1 _9491_/X sky130_fd_sc_hd__mux2_1
X_8442_ _8441_/A _8441_/B _8463_/A vssd1 vssd1 vccd1 vccd1 _8442_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_175_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5654_ _6558_/A vssd1 vssd1 vccd1 vccd1 _8389_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_191_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8373_ _8322_/Y _8373_/B _8373_/C _8373_/D vssd1 vssd1 vccd1 vccd1 _8374_/B sky130_fd_sc_hd__and4b_1
XFILLER_190_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5585_ _5609_/A _5585_/B vssd1 vssd1 vccd1 vccd1 _9709_/D sky130_fd_sc_hd__nor2_1
X_7324_ _7324_/A _7385_/B _7324_/C vssd1 vssd1 vccd1 vccd1 _7324_/X sky130_fd_sc_hd__or3_1
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7255_ _7255_/A _7261_/A vssd1 vssd1 vccd1 vccd1 _7255_/Y sky130_fd_sc_hd__nor2_1
X_6206_ _9576_/Q vssd1 vssd1 vccd1 vccd1 _8001_/A sky130_fd_sc_hd__inv_2
X_7186_ _7186_/A _7192_/A vssd1 vssd1 vccd1 vccd1 _7186_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6137_ _6137_/A vssd1 vssd1 vccd1 vccd1 _6241_/A sky130_fd_sc_hd__clkbuf_4
X_6068_ _6068_/A vssd1 vssd1 vccd1 vccd1 _6068_/Y sky130_fd_sc_hd__inv_2
X_5019_ _5028_/A vssd1 vssd1 vccd1 vccd1 _5019_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9827_ _9929_/CLK _9827_/D vssd1 vssd1 vccd1 vccd1 _9827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9758_ _9909_/CLK _9758_/D vssd1 vssd1 vccd1 vccd1 _9758_/Q sky130_fd_sc_hd__dfxtp_1
X_8709_ _8709_/A _8709_/B vssd1 vssd1 vccd1 vccd1 _8709_/X sky130_fd_sc_hd__or2_1
XFILLER_186_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9689_ _9692_/CLK _9689_/D vssd1 vssd1 vccd1 vccd1 _9689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater86 _9327_/S vssd1 vssd1 vccd1 vccd1 _9291_/S sky130_fd_sc_hd__buf_8
XFILLER_145_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5370_ _5370_/A vssd1 vssd1 vccd1 vccd1 _9725_/D sky130_fd_sc_hd__inv_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7040_ _7015_/X _7034_/X _7015_/X _7034_/X vssd1 vssd1 vccd1 vccd1 _7057_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_clock clock vssd1 vssd1 vccd1 vccd1 clkbuf_0_clock/X sky130_fd_sc_hd__clkbuf_16
X_8991_ _9791_/Q _9908_/Q _9480_/S vssd1 vssd1 vccd1 vccd1 _8991_/X sky130_fd_sc_hd__mux2_1
X_7942_ _9498_/X _7956_/B vssd1 vssd1 vccd1 vccd1 _7942_/Y sky130_fd_sc_hd__nor2_1
X_7873_ _7873_/A _7873_/B vssd1 vssd1 vccd1 vccd1 _7877_/B sky130_fd_sc_hd__or2_1
X_9612_ _9656_/CLK _9612_/D vssd1 vssd1 vccd1 vccd1 _9612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6824_ _6814_/C _6823_/A _6813_/A _6823_/Y vssd1 vssd1 vccd1 vccd1 _6824_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9543_ _9915_/CLK _9543_/D vssd1 vssd1 vccd1 vccd1 _9543_/Q sky130_fd_sc_hd__dfxtp_1
X_6755_ _6755_/A _9095_/X vssd1 vssd1 vccd1 vccd1 _6851_/A sky130_fd_sc_hd__or2_2
XFILLER_23_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9474_ _7095_/X _5808_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9474_/X sky130_fd_sc_hd__mux2_1
X_5706_ input3/X input6/X input7/X input8/X vssd1 vssd1 vccd1 vccd1 _5917_/B sky130_fd_sc_hd__or4_4
X_8425_ _8755_/A _8626_/B _8829_/A _8543_/B vssd1 vssd1 vccd1 vccd1 _8428_/B sky130_fd_sc_hd__o22a_1
XFILLER_163_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6686_ _6682_/X _6685_/X _6682_/X _6685_/X vssd1 vssd1 vccd1 vccd1 _6686_/X sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_1_0_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_clock/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5637_ _9681_/Q vssd1 vssd1 vccd1 vccd1 _8381_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8356_ _7709_/X _9553_/Q _7881_/X _9554_/Q vssd1 vssd1 vccd1 vccd1 _8356_/X sky130_fd_sc_hd__o22a_1
XFILLER_128_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5568_ _5553_/X _5565_/Y _5566_/X _7650_/A _5557_/X vssd1 vssd1 vccd1 vccd1 _5569_/B
+ sky130_fd_sc_hd__o32a_1
X_8287_ _4802_/A _8218_/Y _4798_/A _8217_/X _8286_/X vssd1 vssd1 vccd1 vccd1 _8287_/X
+ sky130_fd_sc_hd__o221a_1
X_7307_ _7303_/A _7303_/B _7372_/B vssd1 vssd1 vccd1 vccd1 _7307_/X sky130_fd_sc_hd__a21o_1
X_7238_ _7247_/A _7238_/B vssd1 vssd1 vccd1 vccd1 _7239_/A sky130_fd_sc_hd__or2_2
X_5499_ _5427_/X _5454_/X _5427_/X _5454_/X vssd1 vssd1 vccd1 vccd1 _5499_/X sky130_fd_sc_hd__a2bb2o_4
X_7169_ _7497_/A _7169_/B vssd1 vssd1 vccd1 vccd1 _7170_/A sky130_fd_sc_hd__or2_4
XFILLER_100_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4870_ _4879_/A vssd1 vssd1 vccd1 vccd1 _4870_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_205_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6540_ _6541_/A _6540_/B vssd1 vssd1 vccd1 vccd1 _6540_/Y sky130_fd_sc_hd__nor2_1
XFILLER_201_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6471_ _9786_/Q _6520_/B _9787_/Q _6521_/B vssd1 vssd1 vccd1 vccd1 _6480_/C sky130_fd_sc_hd__a22o_1
X_8210_ _6416_/A _8209_/Y _6347_/A _8199_/B vssd1 vssd1 vccd1 vccd1 _8210_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9190_ _6532_/Y _9795_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9544_/D sky130_fd_sc_hd__mux2_1
X_5422_ _9365_/X vssd1 vssd1 vccd1 vccd1 _5423_/B sky130_fd_sc_hd__inv_2
XFILLER_160_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8141_ _7810_/A _8119_/Y _8140_/Y vssd1 vssd1 vccd1 vccd1 _8141_/X sky130_fd_sc_hd__a21o_1
X_5353_ _9728_/Q _5353_/B vssd1 vssd1 vccd1 vccd1 _5353_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8072_ _9544_/Q _8072_/B vssd1 vssd1 vccd1 vccd1 _8073_/B sky130_fd_sc_hd__or2_1
XFILLER_87_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5284_ _5279_/B _5271_/X _5283_/Y _5275_/X _5245_/A vssd1 vssd1 vccd1 vccd1 _5285_/A
+ sky130_fd_sc_hd__o32a_1
XINSDIODE2_8 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7023_ _6672_/A _6672_/B _6673_/B vssd1 vssd1 vccd1 vccd1 _7023_/X sky130_fd_sc_hd__a21bo_2
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8974_ _8973_/X _7005_/A _9507_/S vssd1 vssd1 vccd1 vccd1 _8974_/X sky130_fd_sc_hd__mux2_1
X_7925_ _8566_/A vssd1 vssd1 vccd1 vccd1 _8735_/A sky130_fd_sc_hd__buf_2
XFILLER_82_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7856_ _7856_/A _7856_/B vssd1 vssd1 vccd1 vccd1 _7861_/B sky130_fd_sc_hd__or2_1
XPHY_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6807_ _6807_/A _6868_/B _6807_/C vssd1 vssd1 vccd1 vccd1 _6807_/X sky130_fd_sc_hd__or3_1
XFILLER_23_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7787_ _4843_/X _7657_/B _7658_/B vssd1 vssd1 vccd1 vccd1 _7787_/X sky130_fd_sc_hd__a21o_1
X_4999_ _5405_/A vssd1 vssd1 vccd1 vccd1 _5036_/A sky130_fd_sc_hd__buf_2
X_9526_ _9907_/CLK _9526_/D vssd1 vssd1 vccd1 vccd1 _9526_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6738_ _6738_/A _6744_/A vssd1 vssd1 vccd1 vccd1 _6738_/Y sky130_fd_sc_hd__nor2_1
XPHY_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9457_ _8527_/X _8525_/A _9477_/S vssd1 vssd1 vccd1 vccd1 _9457_/X sky130_fd_sc_hd__mux2_2
XFILLER_149_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6669_ _6669_/A vssd1 vssd1 vccd1 vccd1 _6991_/A sky130_fd_sc_hd__inv_2
XFILLER_109_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9388_ _6317_/C _7881_/X _9480_/S vssd1 vssd1 vccd1 vccd1 _9388_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8408_ _9695_/Q _5717_/Y _8384_/Y _8407_/X vssd1 vssd1 vccd1 vccd1 _8408_/X sky130_fd_sc_hd__o22a_1
XFILLER_164_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8339_ _7743_/X _9545_/Q _7723_/X _9546_/Q vssd1 vssd1 vccd1 vccd1 _8339_/X sky130_fd_sc_hd__o22a_1
XFILLER_155_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_16_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _9750_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5971_ _5971_/A vssd1 vssd1 vccd1 vccd1 _5971_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7710_ _4788_/X _6347_/A _7709_/X _6347_/Y vssd1 vssd1 vccd1 vccd1 _7710_/X sky130_fd_sc_hd__o22a_1
X_8690_ _8944_/C _8958_/B _8935_/A _8875_/D vssd1 vssd1 vccd1 vccd1 _8690_/X sky130_fd_sc_hd__o22a_1
X_4922_ _5631_/A vssd1 vssd1 vccd1 vccd1 _4922_/X sky130_fd_sc_hd__clkbuf_4
X_7641_ _7644_/A vssd1 vssd1 vccd1 vccd1 _7648_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4853_ _9896_/Q vssd1 vssd1 vccd1 vccd1 _4853_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4784_ _4799_/A vssd1 vssd1 vccd1 vccd1 _4784_/X sky130_fd_sc_hd__clkbuf_2
X_7572_ _7467_/A _7467_/B _7467_/X vssd1 vssd1 vccd1 vccd1 _7588_/A sky130_fd_sc_hd__a21bo_1
X_9311_ _7886_/Y _9774_/Q _9327_/S vssd1 vssd1 vccd1 vccd1 _9311_/X sky130_fd_sc_hd__mux2_1
X_6523_ _6542_/A vssd1 vssd1 vccd1 vccd1 _6550_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_119_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9242_ _9241_/X _4978_/A _9306_/S vssd1 vssd1 vccd1 vccd1 _9242_/X sky130_fd_sc_hd__mux2_1
X_6454_ _6446_/X _6448_/Y _6451_/Y _6462_/D _6462_/B vssd1 vssd1 vccd1 vccd1 _6454_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_106_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5405_ _5405_/A vssd1 vssd1 vccd1 vccd1 _5910_/A sky130_fd_sc_hd__clkbuf_4
X_9173_ _9172_/X _9781_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9530_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6385_ _9767_/Q _8219_/A vssd1 vssd1 vccd1 vccd1 _8215_/A sky130_fd_sc_hd__or2_2
X_8124_ _8324_/B _8061_/B _8062_/B vssd1 vssd1 vccd1 vccd1 _8124_/X sky130_fd_sc_hd__o21a_1
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5336_ _5336_/A _5346_/A vssd1 vssd1 vccd1 vccd1 _5344_/A sky130_fd_sc_hd__or2_1
X_8055_ _6365_/Y _9530_/Q _4976_/X _8054_/Y vssd1 vssd1 vccd1 vccd1 _8057_/A sky130_fd_sc_hd__a22o_1
X_5267_ _5267_/A vssd1 vssd1 vccd1 vccd1 _5268_/B sky130_fd_sc_hd__inv_2
X_7006_ _7006_/A _7006_/B vssd1 vssd1 vccd1 vccd1 _7006_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5198_ _9759_/Q vssd1 vssd1 vccd1 vccd1 _5198_/X sky130_fd_sc_hd__buf_2
XFILLER_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8957_ _8907_/X _8914_/X _8915_/X _8921_/X vssd1 vssd1 vccd1 vccd1 _8957_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7908_ _8301_/A _7685_/B _9327_/S vssd1 vssd1 vccd1 vccd1 _7908_/X sky130_fd_sc_hd__a21o_1
XFILLER_196_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8888_ _8887_/A _8887_/B _8931_/A vssd1 vssd1 vccd1 vccd1 _8888_/X sky130_fd_sc_hd__a21bo_1
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7839_ _7839_/A vssd1 vssd1 vccd1 vccd1 _7839_/X sky130_fd_sc_hd__buf_4
XPHY_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9509_ _9526_/Q _9008_/X _7930_/Y _9010_/X _8970_/X _9053_/S vssd1 vssd1 vccd1 vccd1
+ _9509_/X sky130_fd_sc_hd__mux4_2
XPHY_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6170_ _6170_/A vssd1 vssd1 vccd1 vccd1 _6171_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5121_ _5138_/A vssd1 vssd1 vccd1 vccd1 _5121_/X sky130_fd_sc_hd__buf_1
XFILLER_111_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5052_ _5069_/A _5052_/B vssd1 vssd1 vccd1 vccd1 _9811_/D sky130_fd_sc_hd__nor2_1
X_9860_ _9930_/CLK _9860_/D vssd1 vssd1 vccd1 vccd1 _9860_/Q sky130_fd_sc_hd__dfxtp_1
X_8811_ _8811_/A _8895_/A vssd1 vssd1 vccd1 vccd1 _8812_/B sky130_fd_sc_hd__or2_1
X_9791_ _9929_/CLK _9791_/D vssd1 vssd1 vccd1 vccd1 _9791_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8742_ _8742_/A vssd1 vssd1 vccd1 vccd1 _8743_/B sky130_fd_sc_hd__inv_2
XFILLER_92_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5954_ _9149_/X _5951_/X _9573_/Q _5952_/X vssd1 vssd1 vccd1 vccd1 _9573_/D sky130_fd_sc_hd__a22o_1
X_8673_ _8546_/A _8629_/A _8776_/A _8766_/B vssd1 vssd1 vccd1 vccd1 _8673_/X sky130_fd_sc_hd__a211o_2
XFILLER_178_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5885_ _5885_/A vssd1 vssd1 vccd1 vccd1 _5885_/X sky130_fd_sc_hd__clkbuf_2
X_4905_ _5631_/A vssd1 vssd1 vccd1 vccd1 _4905_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4836_ _4836_/A vssd1 vssd1 vccd1 vccd1 _4836_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7624_ _7072_/A _7072_/B _7073_/B vssd1 vssd1 vccd1 vccd1 _7624_/X sky130_fd_sc_hd__a21bo_1
XFILLER_166_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7555_ _7527_/X _7528_/X _7529_/X _7554_/Y vssd1 vssd1 vccd1 vccd1 _7555_/Y sky130_fd_sc_hd__o22ai_1
X_4767_ _4799_/A vssd1 vssd1 vccd1 vccd1 _4767_/X sky130_fd_sc_hd__clkbuf_2
X_6506_ _6318_/C _6420_/A _6505_/Y vssd1 vssd1 vccd1 vccd1 _6506_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_174_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7486_ _7209_/X _7485_/Y _7209_/X _7485_/Y vssd1 vssd1 vccd1 vccd1 _7558_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9225_ _9224_/X _7776_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9225_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6437_ _6456_/B vssd1 vssd1 vccd1 vccd1 _6529_/B sky130_fd_sc_hd__inv_2
XFILLER_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6368_ _4976_/X _6364_/Y _6327_/Y _6367_/Y vssd1 vssd1 vccd1 vccd1 _6368_/X sky130_fd_sc_hd__o22a_1
XFILLER_161_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9156_ _6229_/X input24/X _9170_/S vssd1 vssd1 vccd1 vccd1 _9156_/X sky130_fd_sc_hd__mux2_1
X_8107_ _9547_/Q _8075_/B _8076_/B vssd1 vssd1 vccd1 vccd1 _8107_/X sky130_fd_sc_hd__a21bo_1
X_5319_ _9725_/Q vssd1 vssd1 vccd1 vccd1 _5332_/A sky130_fd_sc_hd__inv_2
XFILLER_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6299_ _9594_/Q vssd1 vssd1 vccd1 vccd1 _8046_/A sky130_fd_sc_hd__inv_2
X_9087_ _9086_/X input31/X _9306_/S vssd1 vssd1 vccd1 vccd1 _9087_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8038_ _8038_/A _8044_/B vssd1 vssd1 vccd1 vccd1 _8038_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5670_ _9685_/Q _5658_/X _6571_/A _5662_/X _5660_/X vssd1 vssd1 vccd1 vccd1 _9685_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_187_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7340_ _7334_/A _9475_/X _7313_/C _7389_/B vssd1 vssd1 vccd1 vccd1 _7341_/A sky130_fd_sc_hd__o22a_1
XFILLER_171_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7271_ _7317_/A _9470_/X vssd1 vssd1 vccd1 vccd1 _7277_/C sky130_fd_sc_hd__nor2_1
XFILLER_143_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9010_ _9009_/X _9596_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9010_/X sky130_fd_sc_hd__mux2_1
X_6222_ _8005_/A _6241_/A _8010_/A _6201_/X _6212_/X vssd1 vssd1 vccd1 vccd1 _6222_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_106_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6153_ _6152_/A _6152_/B _6152_/X vssd1 vssd1 vccd1 vccd1 _6153_/Y sky130_fd_sc_hd__a21boi_1
X_5104_ _9799_/Q vssd1 vssd1 vccd1 vccd1 _5104_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6084_ _9859_/Q vssd1 vssd1 vccd1 vccd1 _7990_/A sky130_fd_sc_hd__inv_2
X_5035_ _5035_/A vssd1 vssd1 vccd1 vccd1 _5035_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9912_ _9915_/CLK _9912_/D vssd1 vssd1 vccd1 vccd1 _9912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9843_ _9898_/CLK _9843_/D vssd1 vssd1 vccd1 vccd1 _9843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9774_ _9903_/CLK _9774_/D vssd1 vssd1 vccd1 vccd1 _9774_/Q sky130_fd_sc_hd__dfxtp_1
X_6986_ _6972_/X _6985_/X _6972_/X _6985_/X vssd1 vssd1 vccd1 vccd1 _6986_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8725_ _8958_/A _8725_/B _8725_/C vssd1 vssd1 vccd1 vccd1 _8810_/A sky130_fd_sc_hd__nor3_4
X_5937_ _5937_/A vssd1 vssd1 vccd1 vccd1 _5937_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8656_ _8656_/A vssd1 vssd1 vccd1 vccd1 _8656_/X sky130_fd_sc_hd__buf_2
XFILLER_40_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5868_ _9626_/Q _5865_/X _5026_/X _5866_/X _5867_/X vssd1 vssd1 vccd1 vccd1 _9626_/D
+ sky130_fd_sc_hd__o221a_1
X_7607_ _7604_/A _7604_/B _7604_/X vssd1 vssd1 vccd1 vccd1 _7607_/X sky130_fd_sc_hd__a21bo_1
X_8587_ _8630_/A _8626_/B _8516_/A _8546_/A _8547_/A vssd1 vssd1 vccd1 vccd1 _8628_/A
+ sky130_fd_sc_hd__o32a_1
X_5799_ _9656_/Q _5793_/X _5787_/X _7087_/A _5791_/X vssd1 vssd1 vccd1 vccd1 _9656_/D
+ sky130_fd_sc_hd__o221a_1
X_4819_ _9909_/Q vssd1 vssd1 vccd1 vccd1 _7666_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_181_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7538_ _7476_/X _7537_/X _7476_/X _7537_/X vssd1 vssd1 vccd1 vccd1 _7538_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_162_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7469_ _7459_/X _7460_/X _7461_/X _7468_/X vssd1 vssd1 vccd1 vccd1 _7470_/B sky130_fd_sc_hd__o22ai_4
X_9208_ _9813_/Q _7637_/Y _9528_/Q vssd1 vssd1 vccd1 vccd1 _9208_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput57 _9044_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[12] sky130_fd_sc_hd__clkbuf_2
Xoutput68 _9060_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_88_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput79 _9511_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[3] sky130_fd_sc_hd__clkbuf_2
X_9139_ _9877_/Q _9893_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9139_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6840_ _6785_/A _6785_/B _6786_/B vssd1 vssd1 vccd1 vccd1 _6840_/X sky130_fd_sc_hd__a21bo_1
X_6771_ _6771_/A _6771_/B vssd1 vssd1 vccd1 vccd1 _6782_/A sky130_fd_sc_hd__or2_1
X_8510_ _8510_/A _8531_/B vssd1 vssd1 vccd1 vccd1 _8510_/Y sky130_fd_sc_hd__nor2_1
X_5722_ _9661_/Q vssd1 vssd1 vccd1 vccd1 _5722_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9490_ _8429_/Y _8427_/X _9490_/S vssd1 vssd1 vccd1 vccd1 _9490_/X sky130_fd_sc_hd__mux2_2
X_8441_ _8441_/A _8441_/B vssd1 vssd1 vccd1 vccd1 _8463_/A sky130_fd_sc_hd__nand2_1
X_5653_ _9675_/Q vssd1 vssd1 vccd1 vccd1 _6558_/A sky130_fd_sc_hd__clkbuf_2
X_8372_ _4843_/X _8050_/Y _4847_/X _8052_/Y _8371_/X vssd1 vssd1 vccd1 vccd1 _8373_/D
+ sky130_fd_sc_hd__o221a_1
X_5584_ _5553_/X _5581_/Y _5582_/Y _7647_/A _5577_/X vssd1 vssd1 vccd1 vccd1 _5585_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_175_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7323_ _7323_/A _7323_/B vssd1 vssd1 vccd1 vccd1 _7323_/X sky130_fd_sc_hd__or2_1
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7254_ _7239_/A _7249_/Y _7246_/X _7250_/X vssd1 vssd1 vccd1 vccd1 _7261_/A sky130_fd_sc_hd__o22ai_4
XFILLER_131_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7185_ _7170_/A _7180_/Y _7177_/X _7181_/X vssd1 vssd1 vccd1 vccd1 _7192_/A sky130_fd_sc_hd__o22ai_4
X_6205_ _6221_/A _6204_/Y _6199_/A _6204_/A vssd1 vssd1 vccd1 vccd1 _6205_/X sky130_fd_sc_hd__o22a_1
X_6136_ _6197_/A vssd1 vssd1 vccd1 vccd1 _6137_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6067_ _9857_/Q _6055_/B _6056_/A _6059_/Y vssd1 vssd1 vccd1 vccd1 _6068_/A sky130_fd_sc_hd__o22a_1
X_5018_ _9824_/Q _5011_/X input19/X _5012_/X _5016_/X vssd1 vssd1 vccd1 vccd1 _9824_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_26_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9826_ _9929_/CLK _9826_/D vssd1 vssd1 vccd1 vccd1 _9826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6969_ _6969_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6970_/A sky130_fd_sc_hd__or2_1
X_9757_ _9909_/CLK _9757_/D vssd1 vssd1 vccd1 vccd1 _9757_/Q sky130_fd_sc_hd__dfxtp_2
X_8708_ _8707_/A _8707_/B _8707_/X vssd1 vssd1 vccd1 vccd1 _8708_/X sky130_fd_sc_hd__a21bo_1
XFILLER_167_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9688_ _9692_/CLK _9688_/D vssd1 vssd1 vccd1 vccd1 _9688_/Q sky130_fd_sc_hd__dfxtp_1
X_8639_ _8637_/A _8638_/A _8721_/C _8638_/Y vssd1 vssd1 vccd1 vccd1 _8639_/X sky130_fd_sc_hd__o22a_2
XFILLER_166_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater87 _9331_/S vssd1 vssd1 vccd1 vccd1 _9327_/S sky130_fd_sc_hd__buf_8
XFILLER_157_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8990_ _8989_/X _7005_/A _9507_/S vssd1 vssd1 vccd1 vccd1 _8990_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7941_ _7941_/A _9503_/S vssd1 vssd1 vccd1 vccd1 _7941_/X sky130_fd_sc_hd__or2_1
XFILLER_67_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7872_ _4790_/X _7677_/B _7871_/Y vssd1 vssd1 vccd1 vccd1 _7872_/X sky130_fd_sc_hd__a21o_1
XFILLER_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9611_ _9715_/CLK _9611_/D vssd1 vssd1 vccd1 vccd1 _9611_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6823_ _6823_/A vssd1 vssd1 vccd1 vccd1 _6823_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9542_ _9907_/CLK _9542_/D vssd1 vssd1 vccd1 vccd1 _9542_/Q sky130_fd_sc_hd__dfxtp_1
X_6754_ _6755_/A _9093_/X vssd1 vssd1 vccd1 vccd1 _6760_/C sky130_fd_sc_hd__nor2_2
XFILLER_176_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6685_ _6978_/C _9465_/X _6684_/X vssd1 vssd1 vccd1 vccd1 _6685_/X sky130_fd_sc_hd__or3b_1
X_5705_ _6804_/C _4897_/X _5910_/A _5704_/X vssd1 vssd1 vccd1 vccd1 _9668_/D sky130_fd_sc_hd__o211a_1
X_9473_ _7094_/X _6116_/Y _9475_/S vssd1 vssd1 vccd1 vccd1 _9473_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8424_ _9379_/X vssd1 vssd1 vccd1 vccd1 _8626_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_176_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5636_ _9698_/Q _5631_/X _6982_/A _5635_/X _5632_/X vssd1 vssd1 vccd1 vccd1 _9698_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8355_ _9926_/Q _8092_/Y _7682_/A _8354_/Y vssd1 vssd1 vccd1 vccd1 _8357_/C sky130_fd_sc_hd__a22o_1
XFILLER_117_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5567_ _9712_/Q vssd1 vssd1 vccd1 vccd1 _7650_/A sky130_fd_sc_hd__inv_2
X_5498_ _9403_/X _5497_/X _9403_/X _5497_/X vssd1 vssd1 vccd1 vccd1 _5595_/A sky130_fd_sc_hd__a2bb2oi_1
X_8286_ _9917_/Q _8218_/Y _8285_/Y vssd1 vssd1 vccd1 vccd1 _8286_/X sky130_fd_sc_hd__a21o_1
X_7306_ _7284_/X _7305_/X _7284_/X _7305_/X vssd1 vssd1 vccd1 vccd1 _7306_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_208_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7237_ _7218_/X _7222_/X _7235_/X _7236_/X vssd1 vssd1 vccd1 vccd1 _7237_/X sky130_fd_sc_hd__o22a_1
XFILLER_144_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7168_ _7152_/X _7153_/X _7166_/X _7167_/X vssd1 vssd1 vccd1 vccd1 _7168_/X sky130_fd_sc_hd__o22a_1
X_6119_ _7120_/A vssd1 vssd1 vccd1 vccd1 _6119_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7099_ _7265_/A vssd1 vssd1 vccd1 vccd1 _7491_/A sky130_fd_sc_hd__buf_2
XFILLER_46_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9809_ _9926_/CLK _9809_/D vssd1 vssd1 vccd1 vccd1 _9809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6470_ _6469_/Y _6467_/Y _6374_/B vssd1 vssd1 vccd1 vccd1 _6521_/B sky130_fd_sc_hd__o21a_1
XFILLER_118_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5421_ _9349_/X vssd1 vssd1 vccd1 vccd1 _5423_/A sky130_fd_sc_hd__inv_2
XFILLER_173_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8140_ _7707_/A _8120_/X _8139_/X vssd1 vssd1 vccd1 vccd1 _8140_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5352_ _5352_/A vssd1 vssd1 vccd1 vccd1 _5353_/B sky130_fd_sc_hd__inv_2
XFILLER_114_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8071_ _9543_/Q _8112_/A vssd1 vssd1 vccd1 vccd1 _8072_/B sky130_fd_sc_hd__or2_1
X_5283_ _9740_/Q _5283_/B vssd1 vssd1 vccd1 vccd1 _5283_/Y sky130_fd_sc_hd__nor2_1
X_7022_ _6932_/X _6958_/X _6932_/X _6958_/X vssd1 vssd1 vccd1 vccd1 _7022_/X sky130_fd_sc_hd__a2bb2o_1
XINSDIODE2_9 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8973_ _8972_/X _7490_/A _9506_/S vssd1 vssd1 vccd1 vccd1 _8973_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7924_ _8475_/A vssd1 vssd1 vccd1 vccd1 _8566_/A sky130_fd_sc_hd__buf_1
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7855_ _7673_/A _7673_/B _7854_/Y vssd1 vssd1 vccd1 vccd1 _7855_/X sky130_fd_sc_hd__a21o_1
XPHY_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6806_ _6806_/A _6806_/B vssd1 vssd1 vccd1 vccd1 _6806_/X sky130_fd_sc_hd__or2_1
XFILLER_11_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4998_ _9836_/Q _4994_/X input32/X _4995_/X _4991_/X vssd1 vssd1 vccd1 vccd1 _9836_/D
+ sky130_fd_sc_hd__o221a_1
X_7786_ _4847_/X _7783_/B _7788_/B _7785_/X vssd1 vssd1 vccd1 vccd1 _7786_/X sky130_fd_sc_hd__o211a_1
XPHY_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9525_ _9888_/CLK _9525_/D vssd1 vssd1 vccd1 vccd1 _9525_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6737_ _6722_/A _6732_/Y _6729_/X _6733_/X vssd1 vssd1 vccd1 vccd1 _6744_/A sky130_fd_sc_hd__o22ai_2
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6668_ _6668_/A _6674_/A vssd1 vssd1 vccd1 vccd1 _6668_/Y sky130_fd_sc_hd__nor2_1
X_9456_ _9455_/X _7005_/A _9507_/S vssd1 vssd1 vccd1 vccd1 _9456_/X sky130_fd_sc_hd__mux2_1
X_9387_ _9386_/X _6345_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _9387_/X sky130_fd_sc_hd__mux2_1
X_5619_ _5704_/A _5616_/Y _5617_/Y _7638_/A _5607_/X vssd1 vssd1 vccd1 vccd1 _5620_/B
+ sky130_fd_sc_hd__o32a_1
X_8407_ _9694_/Q _5721_/X _8385_/X _8406_/X vssd1 vssd1 vccd1 vccd1 _8407_/X sky130_fd_sc_hd__o22a_1
X_6599_ _6598_/X _6594_/Y _6982_/A _6982_/B vssd1 vssd1 vccd1 vccd1 _6599_/X sky130_fd_sc_hd__a22o_1
X_8338_ _4798_/X _8102_/Y _4802_/X _8337_/Y vssd1 vssd1 vccd1 vccd1 _8340_/C sky130_fd_sc_hd__a22o_1
XFILLER_136_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8269_ _7726_/A _8244_/Y _8268_/X vssd1 vssd1 vccd1 vccd1 _8269_/X sky130_fd_sc_hd__o21ba_1
XFILLER_171_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5970_ _9518_/Q _5969_/Y _9518_/Q _5969_/Y vssd1 vssd1 vccd1 vccd1 _5971_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4921_ _9867_/Q _4914_/X _9719_/Q _4920_/X _4915_/X vssd1 vssd1 vccd1 vccd1 _9867_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_205_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4852_ _9226_/X _4796_/A _7776_/A _4799_/A _4845_/X vssd1 vssd1 vccd1 vccd1 _9897_/D
+ sky130_fd_sc_hd__o221a_1
X_7640_ _7640_/A _7640_/B vssd1 vssd1 vccd1 vccd1 _7640_/Y sky130_fd_sc_hd__nor2_1
XFILLER_193_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4783_ _9923_/Q vssd1 vssd1 vccd1 vccd1 _7680_/A sky130_fd_sc_hd__clkbuf_2
X_7571_ _7465_/X _7467_/X _7465_/X _7467_/X vssd1 vssd1 vccd1 vccd1 _7587_/A sky130_fd_sc_hd__a2bb2o_1
X_9310_ _9309_/X input33/X _9334_/S vssd1 vssd1 vccd1 vccd1 _9310_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6522_ _6522_/A _6522_/B vssd1 vssd1 vccd1 vccd1 _6522_/Y sky130_fd_sc_hd__nor2_1
X_9241_ _9240_/X _7794_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9241_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6453_ _6453_/A _6453_/B vssd1 vssd1 vccd1 vccd1 _6462_/B sky130_fd_sc_hd__or2_1
XFILLER_9_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9172_ _9844_/Q _6486_/B _9178_/S vssd1 vssd1 vccd1 vccd1 _9172_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5404_ _9716_/Q _5313_/X _5397_/Y _5349_/X vssd1 vssd1 vccd1 vccd1 _9716_/D sky130_fd_sc_hd__o22ai_1
X_8123_ _8123_/A _8123_/B vssd1 vssd1 vccd1 vccd1 _8123_/Y sky130_fd_sc_hd__nand2_1
X_6384_ _9766_/Q _8221_/A vssd1 vssd1 vccd1 vccd1 _8219_/A sky130_fd_sc_hd__or2_1
X_5335_ _5335_/A _5352_/A vssd1 vssd1 vccd1 vccd1 _5346_/A sky130_fd_sc_hd__or2_1
X_8054_ _9530_/Q vssd1 vssd1 vccd1 vccd1 _8054_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5266_ _5266_/A vssd1 vssd1 vccd1 vccd1 _9744_/D sky130_fd_sc_hd__inv_2
XFILLER_141_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7005_ _7005_/A _7005_/B vssd1 vssd1 vccd1 vccd1 _7005_/X sky130_fd_sc_hd__or2_1
XFILLER_87_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5197_ input19/X _5192_/X _6335_/A _5193_/X _5194_/X vssd1 vssd1 vccd1 vccd1 _9760_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8956_ _8954_/X _8955_/Y _8954_/X _8955_/Y vssd1 vssd1 vccd1 vccd1 _8956_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7907_ _4770_/X _7903_/Y _7860_/A _7909_/A vssd1 vssd1 vccd1 vccd1 _7907_/X sky130_fd_sc_hd__o211a_1
XFILLER_83_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8887_ _8887_/A _8887_/B vssd1 vssd1 vccd1 vccd1 _8931_/A sky130_fd_sc_hd__or2_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7838_ _4812_/X _7669_/B _7837_/Y vssd1 vssd1 vccd1 vccd1 _7838_/X sky130_fd_sc_hd__a21o_1
XPHY_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7769_ _7769_/A vssd1 vssd1 vccd1 vccd1 _7769_/Y sky130_fd_sc_hd__inv_2
XPHY_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9508_ _9525_/D _9004_/X _7917_/X _9006_/X _8970_/X _9053_/S vssd1 vssd1 vccd1 vccd1
+ _9508_/X sky130_fd_sc_hd__mux4_2
XPHY_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9439_ _8651_/X _8649_/Y _9477_/S vssd1 vssd1 vccd1 vccd1 _9439_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5120_ _5579_/A _5120_/B vssd1 vssd1 vccd1 vccd1 _9796_/D sky130_fd_sc_hd__nor2_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5051_ _5045_/X _6316_/A _5047_/Y _5050_/X vssd1 vssd1 vccd1 vccd1 _5052_/B sky130_fd_sc_hd__o22a_1
XFILLER_111_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8810_ _8810_/A _8810_/B vssd1 vssd1 vccd1 vccd1 _8895_/A sky130_fd_sc_hd__and2_1
X_9790_ _9929_/CLK _9790_/D vssd1 vssd1 vccd1 vccd1 _9790_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8741_ _8739_/X _8740_/X _8739_/X _8740_/X vssd1 vssd1 vccd1 vccd1 _8742_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5953_ _9150_/X _5951_/X _9574_/Q _5952_/X vssd1 vssd1 vccd1 vccd1 _9574_/D sky130_fd_sc_hd__a22o_1
X_8672_ _8668_/Y _8671_/X _8668_/Y _8671_/X vssd1 vssd1 vccd1 vccd1 _8672_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_178_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5884_ _5884_/A vssd1 vssd1 vccd1 vccd1 _5884_/X sky130_fd_sc_hd__clkbuf_2
X_4904_ _9877_/Q _4897_/X _9729_/Q _4903_/X _4867_/X vssd1 vssd1 vccd1 vccd1 _9877_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4835_ _9903_/Q vssd1 vssd1 vccd1 vccd1 _4835_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7623_ _7596_/A _7596_/B _7597_/B vssd1 vssd1 vccd1 vccd1 _7623_/X sky130_fd_sc_hd__a21bo_1
X_4766_ _4836_/A vssd1 vssd1 vccd1 vccd1 _4799_/A sky130_fd_sc_hd__buf_2
XFILLER_138_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7554_ _7532_/Y _7552_/Y _7553_/Y vssd1 vssd1 vccd1 vccd1 _7554_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6505_ _9800_/Q _6538_/B _6504_/X vssd1 vssd1 vccd1 vccd1 _6505_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_119_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7485_ _7506_/A _7484_/X _7506_/A _7484_/X vssd1 vssd1 vccd1 vccd1 _7485_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9224_ _9748_/Q _9223_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9224_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6436_ _6333_/Y _6435_/Y _8229_/A vssd1 vssd1 vccd1 vccd1 _6456_/B sky130_fd_sc_hd__o21ai_1
X_6367_ _6367_/A vssd1 vssd1 vccd1 vccd1 _6367_/Y sky130_fd_sc_hd__inv_2
X_9155_ _6225_/Y input23/X _9155_/S vssd1 vssd1 vccd1 vccd1 _9155_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8106_ _9548_/Q _8076_/B _8077_/B vssd1 vssd1 vccd1 vccd1 _8106_/X sky130_fd_sc_hd__a21bo_1
XFILLER_88_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5318_ _9726_/Q vssd1 vssd1 vccd1 vccd1 _5333_/A sky130_fd_sc_hd__inv_2
X_6298_ _6295_/X _6297_/X _6295_/X _6297_/X vssd1 vssd1 vccd1 vccd1 _6298_/Y sky130_fd_sc_hd__a2bb2oi_1
X_9086_ _9085_/X _7875_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9086_/X sky130_fd_sc_hd__mux2_1
X_8037_ _9387_/X _8037_/B vssd1 vssd1 vccd1 vccd1 _8037_/Y sky130_fd_sc_hd__nor2_1
X_5249_ _5249_/A _5263_/A vssd1 vssd1 vccd1 vccd1 _5259_/A sky130_fd_sc_hd__or2_2
XFILLER_152_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8939_ _9629_/Q _8908_/Y _5860_/X _8909_/Y _8913_/Y vssd1 vssd1 vccd1 vccd1 _8940_/A
+ sky130_fd_sc_hd__a41o_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_15_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _9708_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7270_ _7268_/X _7269_/X _7268_/X _7269_/X vssd1 vssd1 vccd1 vccd1 _7276_/A sky130_fd_sc_hd__a2bb2o_1
X_6221_ _6221_/A _6221_/B _6221_/C _6221_/D vssd1 vssd1 vccd1 vccd1 _6221_/X sky130_fd_sc_hd__or4_4
X_6152_ _6152_/A _6152_/B vssd1 vssd1 vccd1 vccd1 _6152_/X sky130_fd_sc_hd__or2_2
X_5103_ _5115_/A _5103_/B vssd1 vssd1 vccd1 vccd1 _9800_/D sky130_fd_sc_hd__nor2_1
XFILLER_124_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6083_ _9860_/Q _6081_/Y _7995_/A _9647_/Q vssd1 vssd1 vccd1 vccd1 _6088_/A sky130_fd_sc_hd__a22o_1
X_5034_ _9816_/Q _5028_/X _4978_/X _5030_/X _5024_/X vssd1 vssd1 vccd1 vccd1 _9816_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_111_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9911_ _9915_/CLK _9911_/D vssd1 vssd1 vccd1 vccd1 _9911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9842_ _9898_/CLK _9842_/D vssd1 vssd1 vccd1 vccd1 _9842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9773_ _9903_/CLK _9773_/D vssd1 vssd1 vccd1 vccd1 _9773_/Q sky130_fd_sc_hd__dfxtp_2
X_6985_ _6977_/X _6984_/X _6977_/X _6984_/X vssd1 vssd1 vccd1 vccd1 _6985_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_80_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8724_ _8722_/A _8723_/A _8807_/C _8723_/Y vssd1 vssd1 vccd1 vccd1 _8725_/C sky130_fd_sc_hd__a22o_1
X_5936_ _9161_/X _5930_/X _9585_/Q _5931_/X vssd1 vssd1 vccd1 vccd1 _9585_/D sky130_fd_sc_hd__a22o_1
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8655_ _9632_/Q _8610_/B _8721_/C _8654_/X vssd1 vssd1 vccd1 vccd1 _8655_/X sky130_fd_sc_hd__a31o_1
XFILLER_139_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7606_ _7081_/A _7081_/B _7081_/X vssd1 vssd1 vccd1 vccd1 _7606_/X sky130_fd_sc_hd__a21bo_1
X_5867_ _5891_/A vssd1 vssd1 vccd1 vccd1 _5867_/X sky130_fd_sc_hd__buf_1
XFILLER_193_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8586_ _9631_/Q _8500_/Y _8585_/A _8584_/X _8585_/Y vssd1 vssd1 vccd1 vccd1 _8586_/X
+ sky130_fd_sc_hd__a32o_1
X_4818_ _9079_/X _4809_/X _4816_/X _4810_/X _4817_/X vssd1 vssd1 vccd1 vccd1 _9910_/D
+ sky130_fd_sc_hd__o221a_1
X_5798_ _5798_/A vssd1 vssd1 vccd1 vccd1 _7087_/A sky130_fd_sc_hd__inv_2
X_7537_ _7437_/X _7537_/B vssd1 vssd1 vccd1 vccd1 _7537_/X sky130_fd_sc_hd__and2b_1
X_4749_ input3/X input6/X _5917_/A vssd1 vssd1 vccd1 vccd1 _5815_/D sky130_fd_sc_hd__or3_4
XFILLER_181_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7468_ _7462_/X _7464_/X _7465_/X _7467_/X vssd1 vssd1 vccd1 vccd1 _7468_/X sky130_fd_sc_hd__o22a_1
XFILLER_162_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9207_ _9812_/Q _7636_/Y _9528_/Q vssd1 vssd1 vccd1 vccd1 _9207_/X sky130_fd_sc_hd__mux2_1
X_6419_ _6349_/Y _6418_/Y _8213_/A vssd1 vssd1 vccd1 vccd1 _6420_/A sky130_fd_sc_hd__o21ai_2
XFILLER_107_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput58 _9047_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[13] sky130_fd_sc_hd__clkbuf_2
X_7399_ _7399_/A vssd1 vssd1 vccd1 vccd1 _7400_/C sky130_fd_sc_hd__inv_2
Xoutput69 _9061_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_115_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9138_ _9875_/Q _9891_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9138_/X sky130_fd_sc_hd__mux2_1
X_9069_ _8047_/X _8046_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9069_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6770_ _6759_/A _6759_/B _6759_/X vssd1 vssd1 vccd1 vccd1 _6771_/B sky130_fd_sc_hd__a21bo_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5721_ _5721_/A vssd1 vssd1 vccd1 vccd1 _5721_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8440_ _8440_/A vssd1 vssd1 vccd1 vccd1 _8441_/A sky130_fd_sc_hd__inv_2
X_5652_ _9692_/Q _5645_/X _9676_/Q _5650_/X _5647_/X vssd1 vssd1 vccd1 vccd1 _9692_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8371_ _7778_/B _9529_/Q _4832_/X _8370_/Y vssd1 vssd1 vccd1 vccd1 _8371_/X sky130_fd_sc_hd__o22a_1
X_5583_ _9709_/Q vssd1 vssd1 vccd1 vccd1 _7647_/A sky130_fd_sc_hd__inv_2
XFILLER_175_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7322_ _7324_/C _7320_/X _7576_/A vssd1 vssd1 vccd1 vccd1 _7323_/B sky130_fd_sc_hd__a21oi_1
XFILLER_171_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7253_ _7253_/A vssd1 vssd1 vccd1 vccd1 _7255_/A sky130_fd_sc_hd__inv_2
X_7184_ _7184_/A vssd1 vssd1 vccd1 vccd1 _7186_/A sky130_fd_sc_hd__inv_2
X_6204_ _6204_/A vssd1 vssd1 vccd1 vccd1 _6204_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6135_ _6135_/A vssd1 vssd1 vccd1 vccd1 _6197_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6066_ _6066_/A vssd1 vssd1 vccd1 vccd1 _6066_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5017_ _9825_/Q _5011_/X input20/X _5012_/X _5016_/X vssd1 vssd1 vccd1 vccd1 _9825_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_73_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9825_ _9828_/CLK _9825_/D vssd1 vssd1 vccd1 vccd1 _9825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9756_ _9907_/CLK _9756_/D vssd1 vssd1 vccd1 vccd1 _9756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8707_ _8707_/A _8707_/B vssd1 vssd1 vccd1 vccd1 _8707_/X sky130_fd_sc_hd__or2_1
X_6968_ _6690_/X _6967_/Y _6690_/X _6967_/Y vssd1 vssd1 vccd1 vccd1 _6968_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_53_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9687_ _9699_/CLK _9687_/D vssd1 vssd1 vccd1 vccd1 _9687_/Q sky130_fd_sc_hd__dfxtp_1
X_5919_ _5919_/A _9148_/S vssd1 vssd1 vccd1 vccd1 _5958_/A sky130_fd_sc_hd__or2_4
X_6899_ _6899_/A vssd1 vssd1 vccd1 vccd1 _6925_/A sky130_fd_sc_hd__inv_2
X_8638_ _8638_/A vssd1 vssd1 vccd1 vccd1 _8638_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8569_ _8566_/A _8652_/A _8495_/A _8535_/X _8536_/X vssd1 vssd1 vccd1 vccd1 _8613_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_166_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater88 _9490_/S vssd1 vssd1 vccd1 vccd1 _9477_/S sky130_fd_sc_hd__buf_6
XFILLER_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7940_ _8865_/A vssd1 vssd1 vccd1 vccd1 _8942_/A sky130_fd_sc_hd__buf_4
X_7871_ _7871_/A vssd1 vssd1 vccd1 vccd1 _7871_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6822_ _9614_/Q _6891_/B _6833_/A vssd1 vssd1 vccd1 vccd1 _6823_/A sky130_fd_sc_hd__and3_1
XFILLER_35_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9610_ _9895_/CLK _9610_/D vssd1 vssd1 vccd1 vccd1 _9610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9541_ _9907_/CLK _9541_/D vssd1 vssd1 vccd1 vccd1 _9541_/Q sky130_fd_sc_hd__dfxtp_1
X_6753_ _6751_/X _6752_/X _6751_/X _6752_/X vssd1 vssd1 vccd1 vccd1 _6759_/A sky130_fd_sc_hd__a2bb2o_1
X_6684_ _6982_/D _6981_/B vssd1 vssd1 vccd1 vccd1 _6684_/X sky130_fd_sc_hd__or2_2
X_5704_ _5704_/A _5704_/B _5704_/C vssd1 vssd1 vccd1 vccd1 _5704_/X sky130_fd_sc_hd__or3_1
X_9472_ _7093_/X _5801_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9472_/X sky130_fd_sc_hd__mux2_2
X_8423_ _8605_/A vssd1 vssd1 vccd1 vccd1 _8755_/A sky130_fd_sc_hd__clkbuf_2
X_5635_ _5662_/A vssd1 vssd1 vccd1 vccd1 _5635_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8354_ _9557_/Q vssd1 vssd1 vccd1 vccd1 _8354_/Y sky130_fd_sc_hd__inv_2
X_5566_ _5566_/A _5566_/B vssd1 vssd1 vccd1 vccd1 _5566_/X sky130_fd_sc_hd__and2_1
XFILLER_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8285_ _7856_/A _8220_/X _8284_/X vssd1 vssd1 vccd1 vccd1 _8285_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_104_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7305_ _7299_/A _7294_/X _7298_/Y _7296_/A _7304_/Y vssd1 vssd1 vccd1 vccd1 _7305_/X
+ sky130_fd_sc_hd__o32a_1
X_5497_ _5495_/Y _5496_/Y _5495_/Y _5496_/Y vssd1 vssd1 vccd1 vccd1 _5497_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_208_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7236_ _7218_/X _7222_/X _7218_/X _7222_/X vssd1 vssd1 vccd1 vccd1 _7236_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_86_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7167_ _7152_/X _7153_/X _7152_/X _7153_/X vssd1 vssd1 vccd1 vccd1 _7167_/X sky130_fd_sc_hd__a2bb2o_1
X_6118_ _7089_/A vssd1 vssd1 vccd1 vccd1 _6118_/Y sky130_fd_sc_hd__inv_2
X_7098_ _7331_/A vssd1 vssd1 vccd1 vccd1 _7265_/A sky130_fd_sc_hd__clkbuf_2
X_6049_ _6049_/A vssd1 vssd1 vccd1 vccd1 _6049_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9808_ _9926_/CLK _9808_/D vssd1 vssd1 vccd1 vccd1 _9808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9739_ _9887_/CLK _9739_/D vssd1 vssd1 vccd1 vccd1 _9739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5420_ _9359_/X _9358_/X _9359_/X _9358_/X vssd1 vssd1 vccd1 vccd1 _5420_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5351_ _5351_/A vssd1 vssd1 vccd1 vccd1 _9729_/D sky130_fd_sc_hd__inv_2
XFILLER_160_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8070_ _9542_/Q _8070_/B vssd1 vssd1 vccd1 vccd1 _8112_/A sky130_fd_sc_hd__or2_1
X_5282_ _5282_/A vssd1 vssd1 vccd1 vccd1 _5283_/B sky130_fd_sc_hd__inv_2
XFILLER_99_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7021_ _7019_/X _7020_/X _7019_/X _7020_/X vssd1 vssd1 vccd1 vccd1 _7021_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8972_ _8971_/X _8955_/A _9505_/S vssd1 vssd1 vccd1 vccd1 _8972_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7923_ _9628_/Q vssd1 vssd1 vccd1 vccd1 _8475_/A sky130_fd_sc_hd__inv_2
XFILLER_36_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7854_ _7854_/A vssd1 vssd1 vccd1 vccd1 _7854_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7785_ _7860_/A vssd1 vssd1 vccd1 vccd1 _7785_/X sky130_fd_sc_hd__buf_2
XPHY_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6805_ _6807_/C _6803_/X _7054_/A vssd1 vssd1 vccd1 vccd1 _6806_/B sky130_fd_sc_hd__a21oi_1
XFILLER_63_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4997_ _9837_/Q _4994_/X input33/X _4995_/X _4991_/X vssd1 vssd1 vccd1 vccd1 _9837_/D
+ sky130_fd_sc_hd__o221a_1
X_6736_ _6736_/A vssd1 vssd1 vccd1 vccd1 _6738_/A sky130_fd_sc_hd__inv_2
X_9524_ _9907_/CLK _9524_/D vssd1 vssd1 vccd1 vccd1 _9525_/D sky130_fd_sc_hd__dfxtp_1
XPHY_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6667_ _6652_/A _6662_/Y _6659_/X _6663_/X vssd1 vssd1 vccd1 vccd1 _6674_/A sky130_fd_sc_hd__o22ai_4
XFILLER_109_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9455_ _9454_/X _7490_/A _9506_/S vssd1 vssd1 vccd1 vccd1 _9455_/X sky130_fd_sc_hd__mux2_1
X_9386_ _6317_/B _7885_/X _9480_/S vssd1 vssd1 vccd1 vccd1 _9386_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5618_ _9702_/Q vssd1 vssd1 vccd1 vccd1 _7638_/A sky130_fd_sc_hd__inv_2
X_8406_ _8386_/Y _8405_/Y _9693_/Q _8386_/B vssd1 vssd1 vccd1 vccd1 _8406_/X sky130_fd_sc_hd__a2bb2o_1
X_6598_ _6598_/A vssd1 vssd1 vccd1 vccd1 _6598_/X sky130_fd_sc_hd__buf_1
X_8337_ _9549_/Q vssd1 vssd1 vccd1 vccd1 _8337_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5549_ _5549_/A vssd1 vssd1 vccd1 vccd1 _9350_/S sky130_fd_sc_hd__inv_2
XFILLER_117_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8268_ _7810_/A _8245_/Y _8267_/Y vssd1 vssd1 vccd1 vccd1 _8268_/X sky130_fd_sc_hd__a21bo_1
X_8199_ _8199_/A _8199_/B vssd1 vssd1 vccd1 vccd1 _8200_/B sky130_fd_sc_hd__or2_1
X_7219_ _9471_/X vssd1 vssd1 vccd1 vccd1 _7222_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_100_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4920_ _5662_/A vssd1 vssd1 vccd1 vccd1 _4920_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_52_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4851_ _9897_/Q vssd1 vssd1 vccd1 vccd1 _7776_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4782_ _4796_/A vssd1 vssd1 vccd1 vccd1 _4782_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7570_ _7461_/X _7468_/X _7461_/X _7468_/X vssd1 vssd1 vccd1 vccd1 _7586_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_193_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6521_ _6522_/A _6521_/B vssd1 vssd1 vccd1 vccd1 _6521_/Y sky130_fd_sc_hd__nor2_1
X_9240_ _9752_/Q _9239_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9240_/X sky130_fd_sc_hd__mux2_1
X_6452_ _9791_/Q _6527_/B vssd1 vssd1 vccd1 vccd1 _6462_/D sky130_fd_sc_hd__nand2_1
X_9171_ _6324_/Y _9780_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9529_/D sky130_fd_sc_hd__mux2_1
XFILLER_134_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5403_ _5396_/Y _5349_/X _5313_/X _5402_/X vssd1 vssd1 vccd1 vccd1 _9717_/D sky130_fd_sc_hd__o22ai_1
XFILLER_161_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8122_ _9534_/Q _8062_/B _8063_/B vssd1 vssd1 vccd1 vccd1 _8123_/B sky130_fd_sc_hd__a21boi_2
XFILLER_133_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6383_ _9765_/Q _8223_/A vssd1 vssd1 vccd1 vccd1 _8221_/A sky130_fd_sc_hd__or2_1
X_5334_ _5334_/A _5357_/A vssd1 vssd1 vccd1 vccd1 _5352_/A sky130_fd_sc_hd__or2_1
X_8053_ _8053_/A _9531_/Q vssd1 vssd1 vccd1 vccd1 _8053_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5265_ _5260_/B _5224_/X _5264_/Y _4853_/X _5249_/A vssd1 vssd1 vccd1 vccd1 _5266_/A
+ sky130_fd_sc_hd__o32a_1
X_7004_ _6987_/X _6997_/X _6998_/X _7003_/X vssd1 vssd1 vccd1 vccd1 _7004_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_102_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5196_ _9760_/Q vssd1 vssd1 vccd1 vccd1 _6335_/A sky130_fd_sc_hd__buf_2
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8955_ _8955_/A _8955_/B vssd1 vssd1 vccd1 vccd1 _8955_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7906_ _7906_/A _7906_/B vssd1 vssd1 vccd1 vccd1 _7909_/A sky130_fd_sc_hd__or2_2
X_8886_ _8886_/A vssd1 vssd1 vccd1 vccd1 _8887_/B sky130_fd_sc_hd__inv_2
XFILLER_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7837_ _7837_/A vssd1 vssd1 vccd1 vccd1 _7837_/Y sky130_fd_sc_hd__inv_2
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7768_ _9918_/Q vssd1 vssd1 vccd1 vccd1 _7865_/A sky130_fd_sc_hd__inv_2
XPHY_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7699_ _9924_/Q vssd1 vssd1 vccd1 vccd1 _7891_/A sky130_fd_sc_hd__inv_2
XFILLER_137_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6719_ _6701_/X _6705_/X _6701_/X _6705_/X vssd1 vssd1 vccd1 vccd1 _6719_/X sky130_fd_sc_hd__a2bb2o_1
X_9507_ _9506_/X _9611_/Q _9507_/S vssd1 vssd1 vccd1 vccd1 _9507_/X sky130_fd_sc_hd__mux2_1
XPHY_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9438_ _9437_/X _9775_/Q _9481_/S vssd1 vssd1 vccd1 vccd1 _9438_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9369_ _9368_/X _8955_/A _9505_/S vssd1 vssd1 vccd1 vccd1 _9369_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5050_ _5097_/A vssd1 vssd1 vccd1 vccd1 _5050_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8740_ _8683_/X _8691_/X _8642_/X _8692_/X vssd1 vssd1 vccd1 vccd1 _8740_/X sky130_fd_sc_hd__o22a_1
XFILLER_65_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5952_ _5959_/A vssd1 vssd1 vccd1 vccd1 _5952_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4903_ _5787_/A vssd1 vssd1 vccd1 vccd1 _4903_/X sky130_fd_sc_hd__buf_2
X_8671_ _5843_/X _8500_/Y _8712_/C _8670_/X vssd1 vssd1 vccd1 vccd1 _8671_/X sky130_fd_sc_hd__a31o_1
XFILLER_178_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5883_ _5885_/A vssd1 vssd1 vccd1 vccd1 _5884_/A sky130_fd_sc_hd__inv_2
XFILLER_33_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4834_ _4834_/A vssd1 vssd1 vccd1 vccd1 _4834_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7622_ _7073_/A _7073_/B _7074_/B vssd1 vssd1 vccd1 vccd1 _7622_/X sky130_fd_sc_hd__a21bo_1
XFILLER_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4765_ _4765_/A vssd1 vssd1 vccd1 vccd1 _8301_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_193_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7553_ _7553_/A _7553_/B vssd1 vssd1 vccd1 vccd1 _7553_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6504_ _9800_/Q _6538_/B _6424_/Y _6503_/X vssd1 vssd1 vccd1 vccd1 _6504_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_119_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9223_ _7778_/B _9748_/Q _9327_/S vssd1 vssd1 vccd1 vccd1 _9223_/X sky130_fd_sc_hd__mux2_1
X_7484_ _7263_/X _7482_/X _7217_/X _7483_/X vssd1 vssd1 vccd1 vccd1 _7484_/X sky130_fd_sc_hd__o211a_1
XFILLER_174_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6435_ _6435_/A vssd1 vssd1 vccd1 vccd1 _6435_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6366_ _9845_/Q _6364_/Y _6365_/Y _8184_/B vssd1 vssd1 vccd1 vccd1 _6367_/A sky130_fd_sc_hd__o22a_1
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9154_ _6218_/X input22/X _9155_/S vssd1 vssd1 vccd1 vccd1 _9154_/X sky130_fd_sc_hd__mux2_1
X_9085_ _9771_/Q _9084_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9085_/X sky130_fd_sc_hd__mux2_1
X_8105_ _9549_/Q _8077_/B _8103_/Y vssd1 vssd1 vccd1 vccd1 _8105_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_121_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5317_ _9727_/Q vssd1 vssd1 vccd1 vccd1 _5334_/A sky130_fd_sc_hd__inv_2
XFILLER_0_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6297_ _8040_/A _6193_/A _8042_/A _6142_/A _6296_/X vssd1 vssd1 vccd1 vccd1 _6297_/X
+ sky130_fd_sc_hd__o221a_1
X_8036_ _8036_/A _8044_/B vssd1 vssd1 vccd1 vccd1 _8036_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5248_ _5248_/A _5267_/A vssd1 vssd1 vccd1 vccd1 _5263_/A sky130_fd_sc_hd__or2_1
X_5179_ _5179_/A vssd1 vssd1 vccd1 vccd1 _5179_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8938_ _8938_/A _9422_/X vssd1 vssd1 vccd1 vccd1 _8938_/X sky130_fd_sc_hd__or2_1
XFILLER_56_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8869_ _8867_/X _8868_/X _8867_/X _8868_/X vssd1 vssd1 vccd1 vccd1 _8869_/Y sky130_fd_sc_hd__a2bb2oi_2
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6220_ _9579_/Q _6168_/A _8013_/A _6241_/A vssd1 vssd1 vccd1 vccd1 _6224_/A sky130_fd_sc_hd__a22o_1
XFILLER_131_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6151_ _6125_/Y _6148_/X _7943_/A _6148_/X _6150_/X vssd1 vssd1 vccd1 vccd1 _6152_/B
+ sky130_fd_sc_hd__o221a_1
X_5102_ _5084_/X _6318_/D _5101_/Y _5097_/X vssd1 vssd1 vccd1 vccd1 _5103_/B sky130_fd_sc_hd__o22a_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6082_ _9860_/Q vssd1 vssd1 vccd1 vccd1 _7995_/A sky130_fd_sc_hd__inv_2
X_5033_ _9817_/Q _5028_/X _5032_/X _5030_/X _5024_/X vssd1 vssd1 vccd1 vccd1 _9817_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_111_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9910_ _9910_/CLK _9910_/D vssd1 vssd1 vccd1 vccd1 _9910_/Q sky130_fd_sc_hd__dfxtp_1
X_9841_ _9898_/CLK _9841_/D vssd1 vssd1 vccd1 vccd1 _9841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9772_ _9926_/CLK _9772_/D vssd1 vssd1 vccd1 vccd1 _9772_/Q sky130_fd_sc_hd__dfxtp_1
X_6984_ _6980_/X _6983_/Y _6980_/X _6983_/Y vssd1 vssd1 vccd1 vccd1 _6984_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_80_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8723_ _8723_/A vssd1 vssd1 vccd1 vccd1 _8723_/Y sky130_fd_sc_hd__inv_2
X_5935_ _9162_/X _5930_/X _9586_/Q _5931_/X vssd1 vssd1 vccd1 vccd1 _9586_/D sky130_fd_sc_hd__a22o_1
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8654_ _8875_/A _8773_/D _8807_/A _8725_/B vssd1 vssd1 vccd1 vccd1 _8654_/X sky130_fd_sc_hd__o22a_1
X_5866_ _5866_/A vssd1 vssd1 vccd1 vccd1 _5866_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4817_ _4830_/A vssd1 vssd1 vccd1 vccd1 _4817_/X sky130_fd_sc_hd__clkbuf_2
X_7605_ _7560_/X _7604_/X _7560_/X _7604_/X vssd1 vssd1 vccd1 vccd1 _7605_/Y sky130_fd_sc_hd__a2bb2oi_1
X_8585_ _8585_/A vssd1 vssd1 vccd1 vccd1 _8585_/Y sky130_fd_sc_hd__inv_2
X_5797_ _5736_/X _5747_/X _5736_/X _5747_/X vssd1 vssd1 vccd1 vccd1 _5798_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7536_ _7191_/A _7191_/B _7502_/B vssd1 vssd1 vccd1 vccd1 _7536_/X sky130_fd_sc_hd__a21o_1
X_4748_ _5707_/A _5707_/B _5707_/C input9/X vssd1 vssd1 vccd1 vccd1 _5917_/A sky130_fd_sc_hd__or4_4
XFILLER_174_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7467_ _7467_/A _7467_/B vssd1 vssd1 vccd1 vccd1 _7467_/X sky130_fd_sc_hd__or2_1
X_9206_ _6550_/Y _9811_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9560_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6418_ _6418_/A vssd1 vssd1 vccd1 vccd1 _6418_/Y sky130_fd_sc_hd__inv_2
X_9137_ _9874_/Q _9890_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9137_/X sky130_fd_sc_hd__mux2_1
X_7398_ _7407_/A _7398_/B vssd1 vssd1 vccd1 vccd1 _7399_/A sky130_fd_sc_hd__or2_2
X_6349_ _9769_/Q vssd1 vssd1 vccd1 vccd1 _6349_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput59 _9050_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_88_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9068_ _8045_/Y _8044_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9068_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8019_ _8019_/A _8021_/B vssd1 vssd1 vccd1 vccd1 _8019_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5720_ _9678_/Q vssd1 vssd1 vccd1 vccd1 _5721_/A sky130_fd_sc_hd__inv_2
XFILLER_203_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5651_ _9693_/Q _5645_/X _6576_/A _5650_/X _5647_/X vssd1 vssd1 vccd1 vccd1 _9693_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8370_ _9536_/Q vssd1 vssd1 vccd1 vccd1 _8370_/Y sky130_fd_sc_hd__inv_2
X_5582_ _5582_/A _5582_/B vssd1 vssd1 vccd1 vccd1 _5582_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7321_ _7492_/C _7321_/B _9620_/Q _7321_/D vssd1 vssd1 vccd1 vccd1 _7576_/A sky130_fd_sc_hd__and4_1
X_7252_ _7235_/X _7236_/X _7235_/X _7236_/X vssd1 vssd1 vccd1 vccd1 _7253_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_171_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6203_ _6203_/A _6203_/B vssd1 vssd1 vccd1 vccd1 _6204_/A sky130_fd_sc_hd__nand2_1
X_7183_ _7166_/X _7167_/X _7166_/X _7167_/X vssd1 vssd1 vccd1 vccd1 _7184_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_97_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6134_ _6148_/A vssd1 vssd1 vccd1 vccd1 _6135_/A sky130_fd_sc_hd__buf_1
XFILLER_112_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6065_ _7986_/A _9645_/Q _9858_/Q _6064_/Y vssd1 vssd1 vccd1 vccd1 _6066_/A sky130_fd_sc_hd__o22a_2
X_5016_ _5036_/A vssd1 vssd1 vccd1 vccd1 _5016_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9824_ _9828_/CLK _9824_/D vssd1 vssd1 vccd1 vccd1 _9824_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_14_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _9819_/CLK sky130_fd_sc_hd__clkbuf_16
X_9755_ _9796_/CLK _9755_/D vssd1 vssd1 vccd1 vccd1 _9755_/Q sky130_fd_sc_hd__dfxtp_2
X_6967_ _6995_/A _6966_/X _6995_/A _6966_/X vssd1 vssd1 vccd1 vccd1 _6967_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_14_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8706_ _8619_/A _8621_/Y _8665_/Y _8705_/X vssd1 vssd1 vccd1 vccd1 _8707_/B sky130_fd_sc_hd__a31oi_2
XFILLER_81_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5918_ _5918_/A _7919_/A vssd1 vssd1 vccd1 vccd1 _9148_/S sky130_fd_sc_hd__nor2_8
XFILLER_167_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9686_ _9692_/CLK _9686_/D vssd1 vssd1 vccd1 vccd1 _9686_/Q sky130_fd_sc_hd__dfxtp_1
X_6898_ _6898_/A _6904_/A vssd1 vssd1 vccd1 vccd1 _6898_/Y sky130_fd_sc_hd__nor2_1
XFILLER_194_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8637_ _8637_/A vssd1 vssd1 vccd1 vccd1 _8721_/C sky130_fd_sc_hd__inv_2
X_5849_ _5843_/X _5847_/X _5026_/X _5848_/X _5840_/X vssd1 vssd1 vccd1 vccd1 _9634_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_29_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _9858_/CLK sky130_fd_sc_hd__clkbuf_16
X_8568_ _5860_/X _8656_/A _8566_/X _8567_/Y vssd1 vssd1 vccd1 vccd1 _8568_/X sky130_fd_sc_hd__a31o_1
XFILLER_158_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7519_ _7517_/X _7518_/X _7517_/X _7518_/X vssd1 vssd1 vccd1 vccd1 _7519_/Y sky130_fd_sc_hd__a2bb2oi_1
X_8499_ _8499_/A vssd1 vssd1 vccd1 vccd1 _8499_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater89 _9155_/S vssd1 vssd1 vccd1 vccd1 _9170_/S sky130_fd_sc_hd__buf_8
XFILLER_12_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7870_ _4794_/X _7866_/Y _7860_/X _7873_/B vssd1 vssd1 vccd1 vccd1 _7870_/X sky130_fd_sc_hd__o211a_1
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6821_ _6872_/A _6821_/B vssd1 vssd1 vccd1 vccd1 _6833_/A sky130_fd_sc_hd__or2_1
XFILLER_211_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9540_ _9907_/CLK _9540_/D vssd1 vssd1 vccd1 vccd1 _9540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6752_ _6807_/A _6764_/B vssd1 vssd1 vccd1 vccd1 _6752_/X sky130_fd_sc_hd__or2_1
XFILLER_149_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6683_ _6683_/A vssd1 vssd1 vccd1 vccd1 _6978_/C sky130_fd_sc_hd__buf_2
X_9471_ _7092_/X _5798_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9471_/X sky130_fd_sc_hd__mux2_4
X_5703_ _9848_/Q _5703_/B vssd1 vssd1 vccd1 vccd1 _5704_/C sky130_fd_sc_hd__nor2_2
X_8422_ _8452_/A vssd1 vssd1 vccd1 vccd1 _8605_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5634_ _9682_/Q vssd1 vssd1 vccd1 vccd1 _6982_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8353_ _7885_/X _9555_/Q _7881_/X _9554_/Q vssd1 vssd1 vccd1 vccd1 _8357_/B sky130_fd_sc_hd__a22o_1
XFILLER_191_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5565_ _5565_/A vssd1 vssd1 vccd1 vccd1 _5565_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7304_ _7304_/A _7372_/B vssd1 vssd1 vccd1 vccd1 _7304_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8284_ _7856_/A _8220_/X _8283_/X vssd1 vssd1 vccd1 vccd1 _8284_/X sky130_fd_sc_hd__a21o_1
X_5496_ _5426_/A _5426_/B _5426_/Y vssd1 vssd1 vccd1 vccd1 _5496_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_208_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7235_ _7223_/X _7224_/X _7233_/X _7234_/X vssd1 vssd1 vccd1 vccd1 _7235_/X sky130_fd_sc_hd__o22a_1
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7166_ _7155_/X _7156_/X _7164_/X _7165_/X vssd1 vssd1 vccd1 vccd1 _7166_/X sky130_fd_sc_hd__o22a_1
XFILLER_112_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6117_ _7088_/A vssd1 vssd1 vccd1 vccd1 _6117_/Y sky130_fd_sc_hd__inv_2
X_7097_ _7313_/C vssd1 vssd1 vccd1 vccd1 _7331_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6048_ _6048_/A _6048_/B vssd1 vssd1 vccd1 vccd1 _6049_/A sky130_fd_sc_hd__or2_1
XFILLER_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9807_ _9898_/CLK _9807_/D vssd1 vssd1 vccd1 vccd1 _9807_/Q sky130_fd_sc_hd__dfxtp_1
X_7999_ _7999_/A _8003_/B vssd1 vssd1 vccd1 vccd1 _7999_/X sky130_fd_sc_hd__or2_1
XFILLER_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9738_ _9887_/CLK _9738_/D vssd1 vssd1 vccd1 vccd1 _9738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9669_ _9673_/CLK _9669_/D vssd1 vssd1 vccd1 vccd1 _9669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5350_ _5344_/Y _5313_/X _5347_/Y _5336_/A _5349_/X vssd1 vssd1 vccd1 vccd1 _5351_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5281_ _5281_/A vssd1 vssd1 vccd1 vccd1 _9741_/D sky130_fd_sc_hd__inv_2
XFILLER_141_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7020_ _6673_/A _6673_/B _6991_/B vssd1 vssd1 vccd1 vccd1 _7020_/X sky130_fd_sc_hd__a21o_1
XFILLER_4_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8971_ _7969_/X _6034_/B _9504_/S vssd1 vssd1 vccd1 vccd1 _8971_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7922_ _7922_/A vssd1 vssd1 vccd1 vccd1 _9481_/S sky130_fd_sc_hd__inv_16
XFILLER_67_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7853_ _9915_/Q _7849_/Y _7818_/X _7856_/B vssd1 vssd1 vccd1 vccd1 _7853_/X sky130_fd_sc_hd__o211a_1
XFILLER_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4996_ _9838_/Q _4994_/X input34/X _4995_/X _4991_/X vssd1 vssd1 vccd1 vccd1 _9838_/D
+ sky130_fd_sc_hd__o221a_1
XPHY_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7784_ _7839_/A vssd1 vssd1 vccd1 vccd1 _7860_/A sky130_fd_sc_hd__inv_2
X_6804_ _9611_/Q _6804_/B _6804_/C _9612_/Q vssd1 vssd1 vccd1 vccd1 _7054_/A sky130_fd_sc_hd__and4_1
XFILLER_196_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6735_ _6718_/X _6719_/X _6718_/X _6719_/X vssd1 vssd1 vccd1 vccd1 _6736_/A sky130_fd_sc_hd__a2bb2o_1
X_9523_ _9907_/CLK _9523_/D vssd1 vssd1 vccd1 vccd1 _9523_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9454_ _9453_/X _8955_/A _9505_/S vssd1 vssd1 vccd1 vccd1 _9454_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6666_ _6666_/A vssd1 vssd1 vccd1 vccd1 _6668_/A sky130_fd_sc_hd__inv_2
XFILLER_31_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5617_ _5617_/A _5617_/B vssd1 vssd1 vccd1 vccd1 _5617_/Y sky130_fd_sc_hd__nor2_1
X_9385_ _8696_/X _8694_/A _9490_/S vssd1 vssd1 vccd1 vccd1 _9385_/X sky130_fd_sc_hd__mux2_2
X_8405_ _9692_/Q _6582_/X _8387_/X _8404_/X vssd1 vssd1 vccd1 vccd1 _8405_/Y sky130_fd_sc_hd__o22ai_2
X_6597_ _6596_/Y _6579_/Y _6593_/B vssd1 vssd1 vccd1 vccd1 _6597_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8336_ _7738_/X _9547_/Q _7723_/X _9546_/Q vssd1 vssd1 vccd1 vccd1 _8340_/B sky130_fd_sc_hd__a22o_1
X_5548_ _5548_/A vssd1 vssd1 vccd1 vccd1 _5548_/Y sky130_fd_sc_hd__inv_2
X_8267_ _9905_/Q _8245_/Y _4832_/X _8247_/X _8266_/X vssd1 vssd1 vccd1 vccd1 _8267_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_2_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5479_ _5479_/A vssd1 vssd1 vccd1 vccd1 _5479_/Y sky130_fd_sc_hd__inv_2
X_7218_ _7218_/A _7217_/X vssd1 vssd1 vccd1 vccd1 _7218_/X sky130_fd_sc_hd__or2b_1
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8198_ _6342_/Y _8197_/Y _6397_/A _8199_/B vssd1 vssd1 vccd1 vccd1 _8198_/X sky130_fd_sc_hd__o22a_1
XFILLER_132_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7149_ _9458_/X vssd1 vssd1 vccd1 vccd1 _7494_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_171_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4850_ _9230_/X _4796_/A _7749_/A _4799_/A _4845_/X vssd1 vssd1 vccd1 vccd1 _9898_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4781_ _9318_/X _4763_/X _4780_/X _4767_/X _4778_/X vssd1 vssd1 vccd1 vccd1 _9924_/D
+ sky130_fd_sc_hd__o221a_1
X_6520_ _6522_/A _6520_/B vssd1 vssd1 vccd1 vccd1 _6520_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6451_ _9790_/Q _6526_/B vssd1 vssd1 vccd1 vccd1 _6451_/Y sky130_fd_sc_hd__nor2_1
X_9170_ _6302_/X input40/X _9170_/S vssd1 vssd1 vccd1 vccd1 _9170_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6382_ _9764_/Q _8225_/A vssd1 vssd1 vccd1 vccd1 _8223_/A sky130_fd_sc_hd__or2_1
X_5402_ _9717_/Q _9716_/Q _5396_/Y _5397_/Y vssd1 vssd1 vccd1 vccd1 _5402_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8121_ _9535_/Q _8063_/B _8064_/B vssd1 vssd1 vccd1 vccd1 _8121_/X sky130_fd_sc_hd__a21bo_1
X_5333_ _5333_/A _5361_/A vssd1 vssd1 vccd1 vccd1 _5357_/A sky130_fd_sc_hd__or2_1
XFILLER_114_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8052_ _9531_/Q vssd1 vssd1 vccd1 vccd1 _8052_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5264_ _9744_/Q _5264_/B vssd1 vssd1 vccd1 vccd1 _5264_/Y sky130_fd_sc_hd__nor2_1
X_7003_ _7003_/A _7003_/B vssd1 vssd1 vccd1 vccd1 _7003_/X sky130_fd_sc_hd__or2_1
XFILLER_87_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5195_ input20/X _5192_/X _9761_/Q _5193_/X _5194_/X vssd1 vssd1 vccd1 vccd1 _9761_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8954_ _9633_/Q _8916_/Y _5852_/X _8754_/Y _8920_/Y vssd1 vssd1 vccd1 vccd1 _8954_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_55_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7905_ _7906_/A _7899_/Y _7685_/B vssd1 vssd1 vccd1 vccd1 _7905_/Y sky130_fd_sc_hd__o21ai_1
X_8885_ _8847_/Y _8884_/X _8847_/Y _8884_/X vssd1 vssd1 vccd1 vccd1 _8886_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7836_ _4814_/X _7832_/Y _7818_/X _7840_/B vssd1 vssd1 vccd1 vccd1 _7836_/X sky130_fd_sc_hd__o211a_1
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7767_ _7776_/A _6324_/A _7749_/A _7765_/Y _7766_/Y vssd1 vssd1 vccd1 vccd1 _7772_/C
+ sky130_fd_sc_hd__o221a_1
X_4979_ _9844_/Q _9445_/S _4978_/X _4965_/A _4974_/X vssd1 vssd1 vccd1 vccd1 _9844_/D
+ sky130_fd_sc_hd__o221a_1
XPHY_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6718_ _6706_/X _6707_/X _6716_/X _6717_/X vssd1 vssd1 vccd1 vccd1 _6718_/X sky130_fd_sc_hd__o22a_1
X_7698_ _7831_/A vssd1 vssd1 vccd1 vccd1 _7698_/X sky130_fd_sc_hd__buf_2
X_9506_ _9505_/X _9619_/Q _9506_/S vssd1 vssd1 vccd1 vccd1 _9506_/X sky130_fd_sc_hd__mux2_1
XPHY_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9437_ _9807_/Q _9924_/Q _9480_/S vssd1 vssd1 vccd1 vccd1 _9437_/X sky130_fd_sc_hd__mux2_1
X_6649_ _6631_/X _6632_/X _6631_/X _6632_/X vssd1 vssd1 vccd1 vccd1 _6649_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_109_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9368_ _7974_/X _6041_/Y _9504_/S vssd1 vssd1 vccd1 vccd1 _9368_/X sky130_fd_sc_hd__mux2_1
X_8319_ _7788_/A _9532_/Q _8134_/A _9531_/Q vssd1 vssd1 vccd1 vccd1 _8369_/A sky130_fd_sc_hd__o22a_1
X_9299_ _7868_/Y _9770_/Q _9327_/S vssd1 vssd1 vccd1 vccd1 _9299_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5951_ _5958_/A vssd1 vssd1 vccd1 vccd1 _5951_/X sky130_fd_sc_hd__clkbuf_2
X_8670_ _8773_/A _8584_/B _7967_/A _8625_/B vssd1 vssd1 vccd1 vccd1 _8670_/X sky130_fd_sc_hd__o22a_1
XFILLER_18_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4902_ _9878_/Q _4897_/X _9730_/Q _4900_/X _4867_/X vssd1 vssd1 vccd1 vccd1 _9878_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_52_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5882_ _5882_/A _7914_/A vssd1 vssd1 vccd1 vccd1 _5885_/A sky130_fd_sc_hd__or2_4
XFILLER_33_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4833_ _9254_/X _4822_/X _4832_/X _4824_/X _4830_/X vssd1 vssd1 vccd1 vccd1 _9904_/D
+ sky130_fd_sc_hd__o221a_1
X_7621_ _7597_/A _7597_/B _7598_/B vssd1 vssd1 vccd1 vccd1 _7621_/X sky130_fd_sc_hd__a21bo_1
X_4764_ _9928_/Q vssd1 vssd1 vccd1 vccd1 _4765_/A sky130_fd_sc_hd__buf_2
XFILLER_193_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7552_ _7533_/X _7534_/X _7535_/X _7551_/X vssd1 vssd1 vccd1 vccd1 _7552_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6503_ _5104_/Y _6423_/A _5108_/Y _6428_/A _6502_/Y vssd1 vssd1 vccd1 vccd1 _6503_/X
+ sky130_fd_sc_hd__o221a_1
X_7483_ _7237_/X _7240_/X _7241_/X _7262_/X vssd1 vssd1 vccd1 vccd1 _7483_/X sky130_fd_sc_hd__o22a_1
X_9222_ _9827_/Q _9222_/A1 _9528_/Q vssd1 vssd1 vccd1 vccd1 _9222_/X sky130_fd_sc_hd__mux2_1
X_6434_ _9794_/Q _6531_/B vssd1 vssd1 vccd1 vccd1 _6465_/C sky130_fd_sc_hd__or2_1
XFILLER_146_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6365_ _9845_/Q vssd1 vssd1 vccd1 vccd1 _6365_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9153_ _6214_/Y input21/X _9155_/S vssd1 vssd1 vccd1 vccd1 _9153_/X sky130_fd_sc_hd__mux2_1
X_6296_ _6296_/A _6296_/B vssd1 vssd1 vccd1 vccd1 _6296_/X sky130_fd_sc_hd__or2_1
X_9084_ _7872_/X _9771_/Q _9327_/S vssd1 vssd1 vccd1 vccd1 _9084_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8104_ _8102_/Y _8103_/Y _8079_/B vssd1 vssd1 vccd1 vccd1 _8104_/X sky130_fd_sc_hd__o21a_1
XFILLER_88_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5316_ _9728_/Q vssd1 vssd1 vccd1 vccd1 _5335_/A sky130_fd_sc_hd__inv_2
X_8035_ _8046_/B vssd1 vssd1 vccd1 vccd1 _8044_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_88_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5247_ _5247_/A _5272_/A vssd1 vssd1 vccd1 vccd1 _5267_/A sky130_fd_sc_hd__or2_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5178_ _5178_/A vssd1 vssd1 vccd1 vccd1 _5178_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8937_ _8933_/X _8936_/X _8933_/X _8936_/X vssd1 vssd1 vccd1 vccd1 _8937_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8868_ _8734_/X _8827_/A _8829_/A _8959_/B vssd1 vssd1 vccd1 vccd1 _8868_/X sky130_fd_sc_hd__a211o_1
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8799_ _8767_/X _8770_/X _8771_/X _8783_/X vssd1 vssd1 vccd1 vccd1 _8799_/X sky130_fd_sc_hd__o22a_1
X_7819_ _7819_/A _7819_/B vssd1 vssd1 vccd1 vccd1 _7823_/B sky130_fd_sc_hd__or2_2
XFILLER_12_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6150_ _6150_/A _6150_/B vssd1 vssd1 vccd1 vccd1 _6150_/X sky130_fd_sc_hd__or2_1
X_5101_ _9832_/Q vssd1 vssd1 vccd1 vccd1 _5101_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6081_ _9647_/Q vssd1 vssd1 vccd1 vccd1 _6081_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5032_ _5032_/A vssd1 vssd1 vccd1 vccd1 _5032_/X sky130_fd_sc_hd__buf_4
X_9840_ _9898_/CLK _9840_/D vssd1 vssd1 vccd1 vccd1 _9840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9771_ _9903_/CLK _9771_/D vssd1 vssd1 vccd1 vccd1 _9771_/Q sky130_fd_sc_hd__dfxtp_2
X_6983_ _6981_/Y _6982_/X _6981_/Y _6982_/X vssd1 vssd1 vccd1 vccd1 _6983_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8722_ _8722_/A vssd1 vssd1 vccd1 vccd1 _8807_/C sky130_fd_sc_hd__inv_2
X_5934_ _9163_/X _5930_/X _9587_/Q _5931_/X vssd1 vssd1 vccd1 vccd1 _9587_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8653_ _8773_/B vssd1 vssd1 vccd1 vccd1 _8725_/B sky130_fd_sc_hd__buf_2
XFILLER_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5865_ _5865_/A vssd1 vssd1 vccd1 vccd1 _5865_/X sky130_fd_sc_hd__clkbuf_2
X_4816_ _9910_/Q vssd1 vssd1 vccd1 vccd1 _4816_/X sky130_fd_sc_hd__clkbuf_2
X_7604_ _7604_/A _7604_/B vssd1 vssd1 vccd1 vccd1 _7604_/X sky130_fd_sc_hd__or2_1
X_8584_ _8606_/A _8584_/B vssd1 vssd1 vccd1 vccd1 _8584_/X sky130_fd_sc_hd__or2_1
X_5796_ _9657_/Q _5793_/X _5787_/X _7088_/A _5791_/X vssd1 vssd1 vccd1 vccd1 _9657_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_147_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4747_ input8/X vssd1 vssd1 vccd1 vccd1 _5815_/B sky130_fd_sc_hd__inv_2
X_7535_ _7533_/X _7534_/X _7533_/X _7534_/X vssd1 vssd1 vccd1 vccd1 _7535_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7466_ _7367_/A _7367_/B _7367_/X vssd1 vssd1 vccd1 vccd1 _7467_/B sky130_fd_sc_hd__a21bo_1
X_9205_ _6549_/Y _9810_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9559_/D sky130_fd_sc_hd__mux2_1
X_6417_ _9770_/Q _8213_/A _6414_/Y vssd1 vssd1 vccd1 vccd1 _6540_/B sky130_fd_sc_hd__a21oi_4
XFILLER_134_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7397_ _7382_/X _7384_/X _7395_/X _7396_/X vssd1 vssd1 vccd1 vccd1 _7397_/X sky130_fd_sc_hd__o22a_1
XFILLER_162_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6348_ _9770_/Q vssd1 vssd1 vccd1 vccd1 _6348_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9136_ _9873_/Q _9889_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9136_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9067_ _8043_/Y _8042_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9067_/X sky130_fd_sc_hd__mux2_1
X_6279_ _9590_/Q vssd1 vssd1 vccd1 vccd1 _8038_/A sky130_fd_sc_hd__inv_2
X_8018_ _9434_/X _8022_/B vssd1 vssd1 vccd1 vccd1 _8018_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5650_ _5662_/A vssd1 vssd1 vccd1 vccd1 _5650_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_203_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5581_ _5581_/A vssd1 vssd1 vccd1 vccd1 _5581_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7320_ _7314_/A _7334_/B _9620_/Q _7408_/B vssd1 vssd1 vccd1 vccd1 _7320_/X sky130_fd_sc_hd__o211a_1
XFILLER_116_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7251_ _7246_/X _7250_/X _7246_/X _7250_/X vssd1 vssd1 vccd1 vccd1 _7428_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_171_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6202_ _7988_/A _6201_/X _7993_/A _6201_/X _6189_/B vssd1 vssd1 vccd1 vccd1 _6203_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_131_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7182_ _7177_/X _7181_/X _7177_/X _7181_/X vssd1 vssd1 vccd1 vccd1 _7503_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_112_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6133_ _9566_/Q _6146_/A _7943_/A _6148_/A vssd1 vssd1 vccd1 vccd1 _6150_/B sky130_fd_sc_hd__a22o_1
XFILLER_97_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6064_ _9645_/Q vssd1 vssd1 vccd1 vccd1 _6064_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5015_ _9826_/Q _5011_/X input21/X _5012_/X _5008_/X vssd1 vssd1 vccd1 vccd1 _9826_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_97_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9823_ _9929_/CLK _9823_/D vssd1 vssd1 vccd1 vccd1 _9823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9754_ _9907_/CLK _9754_/D vssd1 vssd1 vccd1 vccd1 _9754_/Q sky130_fd_sc_hd__dfxtp_1
X_6966_ _6746_/X _6964_/X _6700_/X _6965_/X vssd1 vssd1 vccd1 vccd1 _6966_/X sky130_fd_sc_hd__o211a_1
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8705_ _8619_/B _8663_/Y _8662_/Y vssd1 vssd1 vccd1 vccd1 _8705_/X sky130_fd_sc_hd__o21a_1
XFILLER_179_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5917_ _5917_/A _5917_/B _7918_/A vssd1 vssd1 vccd1 vccd1 _7919_/A sky130_fd_sc_hd__or3_4
XFILLER_194_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9685_ _9692_/CLK _9685_/D vssd1 vssd1 vccd1 vccd1 _9685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6897_ _6882_/A _6892_/Y _6889_/X _6893_/X vssd1 vssd1 vccd1 vccd1 _6904_/A sky130_fd_sc_hd__o22ai_4
XFILLER_194_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8636_ _8624_/X _8635_/X _8624_/X _8635_/X vssd1 vssd1 vccd1 vccd1 _8638_/A sky130_fd_sc_hd__a2bb2o_1
X_5848_ _5848_/A vssd1 vssd1 vccd1 vccd1 _5848_/X sky130_fd_sc_hd__buf_1
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8567_ _5860_/X _8656_/A _8566_/X vssd1 vssd1 vccd1 vccd1 _8567_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_166_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5779_ _5779_/A vssd1 vssd1 vccd1 vccd1 _7109_/A sky130_fd_sc_hd__inv_2
XFILLER_21_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7518_ _7518_/A _9415_/X vssd1 vssd1 vccd1 vccd1 _7518_/X sky130_fd_sc_hd__or2_1
X_8498_ _5858_/X _8610_/B _8536_/C _8497_/X vssd1 vssd1 vccd1 vccd1 _8498_/X sky130_fd_sc_hd__a31o_1
XFILLER_135_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7449_ _7446_/X _7447_/X _7446_/X _7447_/X vssd1 vssd1 vccd1 vccd1 _7449_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_174_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9119_ _9603_/Q input46/X _9667_/Q vssd1 vssd1 vccd1 vccd1 _9119_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6820_ _6806_/X _6807_/X _6806_/X _6807_/X vssd1 vssd1 vccd1 vccd1 _6820_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_35_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6751_ _6755_/A _9092_/X vssd1 vssd1 vccd1 vccd1 _6751_/X sky130_fd_sc_hd__or2_1
XFILLER_35_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6682_ _6682_/A _6681_/X vssd1 vssd1 vccd1 vccd1 _6682_/X sky130_fd_sc_hd__or2b_1
X_9470_ _7091_/X _6117_/Y _9475_/S vssd1 vssd1 vccd1 vccd1 _9470_/X sky130_fd_sc_hd__mux2_4
X_5702_ _9635_/Q vssd1 vssd1 vccd1 vccd1 _5703_/B sky130_fd_sc_hd__inv_2
X_8421_ _8469_/B _8580_/B _9628_/Q _9627_/Q vssd1 vssd1 vccd1 vccd1 _8426_/A sky130_fd_sc_hd__and4b_1
XFILLER_176_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5633_ _9699_/Q _5631_/X _9683_/Q _4920_/X _5632_/X vssd1 vssd1 vccd1 vccd1 _9699_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8352_ _4765_/A _8088_/Y _7684_/A _8048_/Y vssd1 vssd1 vccd1 vccd1 _8357_/A sky130_fd_sc_hd__a22o_1
X_5564_ _5579_/A _5564_/B vssd1 vssd1 vccd1 vccd1 _9713_/D sky130_fd_sc_hd__nor2_1
XFILLER_163_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7303_ _7303_/A _7303_/B vssd1 vssd1 vccd1 vccd1 _7372_/B sky130_fd_sc_hd__nor2_2
XFILLER_208_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8283_ _7738_/A _8222_/X _8282_/Y vssd1 vssd1 vccd1 vccd1 _8283_/X sky130_fd_sc_hd__a21bo_1
X_5495_ _5495_/A vssd1 vssd1 vccd1 vccd1 _5495_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7234_ _7234_/A _7283_/B _7234_/C vssd1 vssd1 vccd1 vccd1 _7234_/X sky130_fd_sc_hd__or3_1
XFILLER_144_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7165_ _7487_/C _7494_/B _7165_/C vssd1 vssd1 vccd1 vccd1 _7165_/X sky130_fd_sc_hd__or3_1
XFILLER_100_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6116_ _7085_/A vssd1 vssd1 vccd1 vccd1 _6116_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7096_ _9622_/Q vssd1 vssd1 vccd1 vccd1 _7313_/C sky130_fd_sc_hd__inv_2
X_6047_ _6047_/A vssd1 vssd1 vccd1 vccd1 _6048_/B sky130_fd_sc_hd__inv_2
XFILLER_85_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9806_ _9836_/CLK _9806_/D vssd1 vssd1 vccd1 vccd1 _9806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7998_ _9450_/X _8002_/B vssd1 vssd1 vccd1 vccd1 _7998_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9737_ _9887_/CLK _9737_/D vssd1 vssd1 vccd1 vccd1 _9737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6949_ _6946_/X _6948_/X _6946_/X _6948_/X vssd1 vssd1 vccd1 vccd1 _6949_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_179_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9668_ _9715_/CLK _9668_/D vssd1 vssd1 vccd1 vccd1 _9668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8619_ _8619_/A _8619_/B vssd1 vssd1 vccd1 vccd1 _8620_/A sky130_fd_sc_hd__or2_1
XFILLER_194_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9599_ _9895_/CLK _9599_/D vssd1 vssd1 vccd1 vccd1 _9599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _9929_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5280_ _5273_/B _5271_/X _5279_/Y _5275_/X _5246_/A vssd1 vssd1 vccd1 vccd1 _5281_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_141_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8970_ _8030_/B _9052_/S _9053_/S vssd1 vssd1 vccd1 vccd1 _8970_/X sky130_fd_sc_hd__mux2_8
XFILLER_67_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _9879_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7921_ _7921_/A vssd1 vssd1 vccd1 vccd1 _9052_/S sky130_fd_sc_hd__buf_4
XFILLER_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7852_ _7852_/A _7852_/B vssd1 vssd1 vccd1 vccd1 _7856_/B sky130_fd_sc_hd__or2_2
XFILLER_63_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4995_ _5004_/A vssd1 vssd1 vccd1 vccd1 _4995_/X sky130_fd_sc_hd__clkbuf_2
X_7783_ _9899_/Q _7783_/B vssd1 vssd1 vccd1 vccd1 _7788_/B sky130_fd_sc_hd__nand2_2
X_6803_ _6796_/C _6800_/A _9612_/Q _6891_/B vssd1 vssd1 vccd1 vccd1 _6803_/X sky130_fd_sc_hd__o211a_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9522_ _9930_/CLK _9522_/D vssd1 vssd1 vccd1 vccd1 _9522_/Q sky130_fd_sc_hd__dfxtp_1
X_6734_ _6729_/X _6733_/X _6729_/X _6733_/X vssd1 vssd1 vccd1 vccd1 _6911_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9453_ _7995_/X _6081_/Y _9504_/S vssd1 vssd1 vccd1 vccd1 _9453_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8404_ _9691_/Q _6551_/Y _8389_/Y _8403_/X vssd1 vssd1 vccd1 vccd1 _8404_/X sky130_fd_sc_hd__o22a_1
X_6665_ _6648_/X _6649_/X _6648_/X _6649_/X vssd1 vssd1 vccd1 vccd1 _6666_/A sky130_fd_sc_hd__a2bb2o_1
X_5616_ _5616_/A vssd1 vssd1 vccd1 vccd1 _5616_/Y sky130_fd_sc_hd__inv_2
X_9384_ _8842_/X _8840_/A _9490_/S vssd1 vssd1 vccd1 vccd1 _9384_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6596_ _6596_/A vssd1 vssd1 vccd1 vccd1 _6596_/Y sky130_fd_sc_hd__inv_2
X_8335_ _4790_/X _8333_/Y _4794_/X _8334_/Y vssd1 vssd1 vccd1 vccd1 _8340_/A sky130_fd_sc_hd__a22o_1
X_5547_ _9423_/X _5546_/Y _9423_/X _5546_/Y vssd1 vssd1 vccd1 vccd1 _5548_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8266_ _4835_/X _8248_/Y _9904_/Q _8247_/X _8265_/X vssd1 vssd1 vccd1 vccd1 _8266_/X
+ sky130_fd_sc_hd__a221o_1
X_5478_ _9384_/X _5477_/X _9384_/X _5477_/X vssd1 vssd1 vccd1 vccd1 _5566_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7217_ _7522_/A _7283_/B _7490_/A _7238_/B vssd1 vssd1 vccd1 vccd1 _7217_/X sky130_fd_sc_hd__or4_4
X_8197_ _8197_/A _8199_/B vssd1 vssd1 vccd1 vccd1 _8197_/Y sky130_fd_sc_hd__nor2_1
XFILLER_132_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7148_ _9625_/Q _7135_/Y _5872_/X _7137_/Y _7147_/Y vssd1 vssd1 vccd1 vccd1 _7148_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_48_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7079_ _7079_/A _7079_/B vssd1 vssd1 vccd1 vccd1 _7080_/B sky130_fd_sc_hd__or2_1
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4780_ _9924_/Q vssd1 vssd1 vccd1 vccd1 _4780_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6450_ _6453_/B vssd1 vssd1 vccd1 vccd1 _6526_/B sky130_fd_sc_hd__inv_2
X_6381_ _9763_/Q _8227_/A vssd1 vssd1 vccd1 vccd1 _8225_/A sky130_fd_sc_hd__or2_2
X_5401_ _5401_/A vssd1 vssd1 vccd1 vccd1 _9718_/D sky130_fd_sc_hd__inv_2
XFILLER_133_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8120_ _9536_/Q _8064_/B _8065_/B vssd1 vssd1 vccd1 vccd1 _8120_/X sky130_fd_sc_hd__a21bo_1
X_5332_ _5332_/A _5367_/A vssd1 vssd1 vccd1 vccd1 _5361_/A sky130_fd_sc_hd__or2_1
XFILLER_154_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8051_ _8051_/A _9532_/Q vssd1 vssd1 vccd1 vccd1 _8051_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5263_ _5263_/A vssd1 vssd1 vccd1 vccd1 _5264_/B sky130_fd_sc_hd__inv_2
XFILLER_205_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7002_ _6684_/X _7000_/X _6620_/A _7001_/X vssd1 vssd1 vccd1 vccd1 _7003_/B sky130_fd_sc_hd__o22a_1
X_5194_ _5206_/A vssd1 vssd1 vccd1 vccd1 _5194_/X sky130_fd_sc_hd__buf_1
XFILLER_68_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8953_ _5843_/X _8656_/X _8893_/C _8952_/Y vssd1 vssd1 vccd1 vccd1 _8953_/X sky130_fd_sc_hd__a31o_1
X_7904_ _7902_/A _7902_/B _7790_/X _7903_/Y vssd1 vssd1 vccd1 vccd1 _7904_/Y sky130_fd_sc_hd__a211oi_4
X_8884_ _8927_/A _8927_/B _8883_/Y vssd1 vssd1 vccd1 vccd1 _8884_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7835_ _7835_/A _7835_/B vssd1 vssd1 vccd1 vccd1 _7840_/B sky130_fd_sc_hd__or2_2
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7766_ _4835_/X _7748_/Y _7891_/A _5162_/X vssd1 vssd1 vccd1 vccd1 _7766_/Y sky130_fd_sc_hd__a22oi_1
X_4978_ _4978_/A vssd1 vssd1 vccd1 vccd1 _4978_/X sky130_fd_sc_hd__clkbuf_4
X_9505_ _9504_/X _9627_/Q _9505_/S vssd1 vssd1 vccd1 vccd1 _9505_/X sky130_fd_sc_hd__mux2_1
XPHY_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6717_ _7006_/A _6766_/B _6717_/C vssd1 vssd1 vccd1 vccd1 _6717_/X sky130_fd_sc_hd__or3_1
X_7697_ _9910_/Q vssd1 vssd1 vccd1 vccd1 _7831_/A sky130_fd_sc_hd__inv_2
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9436_ _9435_/X _6350_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _9436_/X sky130_fd_sc_hd__mux2_1
X_6648_ _6634_/X _6637_/X _6646_/X _6647_/X vssd1 vssd1 vccd1 vccd1 _6648_/X sky130_fd_sc_hd__o22a_1
X_9367_ _9366_/X _6339_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _9367_/X sky130_fd_sc_hd__mux2_2
XFILLER_152_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8318_ _7797_/A _9534_/Q _7793_/A _9533_/Q vssd1 vssd1 vccd1 vccd1 _8369_/C sky130_fd_sc_hd__o22a_1
X_6579_ _6592_/B vssd1 vssd1 vccd1 vccd1 _6579_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9298_ _9297_/X input29/X _9306_/S vssd1 vssd1 vccd1 vccd1 _9298_/X sky130_fd_sc_hd__mux2_1
X_8249_ _6371_/A _8209_/Y _8236_/B vssd1 vssd1 vccd1 vccd1 _8249_/X sky130_fd_sc_hd__o21a_1
XFILLER_105_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5950_ _9151_/X _5944_/X _9575_/Q _5945_/X vssd1 vssd1 vccd1 vccd1 _9575_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4901_ _9879_/Q _4897_/X _9731_/Q _4900_/X _4867_/X vssd1 vssd1 vccd1 vccd1 _9879_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7620_ _7074_/A _7074_/B _7075_/B vssd1 vssd1 vccd1 vccd1 _7620_/X sky130_fd_sc_hd__a21bo_1
X_5881_ _5881_/A _5917_/B vssd1 vssd1 vccd1 vccd1 _7914_/A sky130_fd_sc_hd__or2_4
X_4832_ _9904_/Q vssd1 vssd1 vccd1 vccd1 _4832_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4763_ _4796_/A vssd1 vssd1 vccd1 vccd1 _4763_/X sky130_fd_sc_hd__clkbuf_2
X_7551_ _7536_/X _7538_/X _7539_/X _7550_/X vssd1 vssd1 vccd1 vccd1 _7551_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6502_ _9797_/Q _6534_/B _9798_/Q _6535_/B _6501_/Y vssd1 vssd1 vccd1 vccd1 _6502_/Y
+ sky130_fd_sc_hd__o221ai_2
X_7482_ _7482_/A _7482_/B vssd1 vssd1 vccd1 vccd1 _7482_/X sky130_fd_sc_hd__or2_1
X_9221_ _9826_/Q _7652_/Y _9528_/Q vssd1 vssd1 vccd1 vccd1 _9221_/X sky130_fd_sc_hd__mux2_1
X_6433_ _6331_/A _8229_/A _6430_/Y vssd1 vssd1 vccd1 vccd1 _6531_/B sky130_fd_sc_hd__a21oi_2
XFILLER_161_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6364_ _9750_/Q vssd1 vssd1 vccd1 vccd1 _6364_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9152_ _6209_/X input20/X _9155_/S vssd1 vssd1 vccd1 vccd1 _9152_/X sky130_fd_sc_hd__mux2_1
X_6295_ _9593_/Q _6171_/A _8044_/A _6193_/A vssd1 vssd1 vccd1 vccd1 _6295_/X sky130_fd_sc_hd__a22o_1
X_8103_ _8103_/A vssd1 vssd1 vccd1 vccd1 _8103_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9083_ _9082_/X input24/X _9294_/S vssd1 vssd1 vccd1 vccd1 _9083_/X sky130_fd_sc_hd__mux2_1
X_5315_ _9729_/Q vssd1 vssd1 vccd1 vccd1 _5336_/A sky130_fd_sc_hd__inv_2
X_8034_ _9389_/X _8037_/B vssd1 vssd1 vccd1 vccd1 _8034_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5246_ _5246_/A _5278_/A vssd1 vssd1 vccd1 vccd1 _5272_/A sky130_fd_sc_hd__or2_1
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5177_ _9768_/Q vssd1 vssd1 vccd1 vccd1 _6350_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8936_ _8934_/Y _8935_/X _8934_/Y _8935_/X vssd1 vssd1 vccd1 vccd1 _8936_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8867_ _8751_/X _8866_/X _8751_/X _8866_/X vssd1 vssd1 vccd1 vccd1 _8867_/X sky130_fd_sc_hd__a2bb2o_2
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8798_ _8797_/A _8797_/B _8845_/A vssd1 vssd1 vccd1 vccd1 _8798_/X sky130_fd_sc_hd__a21o_1
X_7818_ _7860_/A vssd1 vssd1 vccd1 vccd1 _7818_/X sky130_fd_sc_hd__buf_2
XFILLER_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7749_ _7749_/A vssd1 vssd1 vccd1 vccd1 _8322_/A sky130_fd_sc_hd__inv_2
XFILLER_101_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9419_ _8891_/X _8890_/A _9477_/S vssd1 vssd1 vccd1 vccd1 _9419_/X sky130_fd_sc_hd__mux2_2
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5100_ _9800_/Q vssd1 vssd1 vccd1 vccd1 _6318_/D sky130_fd_sc_hd__inv_2
XFILLER_124_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6080_ _6076_/Y _6079_/X _6076_/Y _6079_/X vssd1 vssd1 vccd1 vccd1 _6080_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5031_ _9818_/Q _5028_/X _5029_/X _5030_/X _5024_/X vssd1 vssd1 vccd1 vccd1 _9818_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_111_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9770_ _9917_/CLK _9770_/D vssd1 vssd1 vccd1 vccd1 _9770_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_65_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8721_ _8776_/A _8773_/D _8721_/C vssd1 vssd1 vccd1 vccd1 _8723_/A sky130_fd_sc_hd__or3_4
X_6982_ _6982_/A _6982_/B _6982_/C _6982_/D vssd1 vssd1 vccd1 vccd1 _6982_/X sky130_fd_sc_hd__or4_4
XFILLER_202_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5933_ _9164_/X _5930_/X _9588_/Q _5931_/X vssd1 vssd1 vccd1 vccd1 _9588_/D sky130_fd_sc_hd__a22o_1
XFILLER_202_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8652_ _8652_/A vssd1 vssd1 vccd1 vccd1 _8773_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_178_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5864_ _5866_/A vssd1 vssd1 vccd1 vccd1 _5865_/A sky130_fd_sc_hd__inv_2
X_8583_ _8630_/A _8625_/B vssd1 vssd1 vccd1 vccd1 _8585_/A sky130_fd_sc_hd__or2_1
XFILLER_178_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4815_ _9278_/X _4809_/X _4814_/X _4810_/X _4806_/X vssd1 vssd1 vccd1 vccd1 _9911_/D
+ sky130_fd_sc_hd__o221a_1
X_7603_ _7603_/A _7603_/B vssd1 vssd1 vccd1 vccd1 _7604_/B sky130_fd_sc_hd__or2_1
X_5795_ _5748_/X _5794_/X _5748_/X _5794_/X vssd1 vssd1 vccd1 vccd1 _7088_/A sky130_fd_sc_hd__o2bb2a_2
X_7534_ _7145_/A _7512_/X _7145_/A _7512_/X vssd1 vssd1 vccd1 vccd1 _7534_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_119_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4746_ input5/X input4/X _4856_/C _4929_/C vssd1 vssd1 vccd1 vccd1 _5147_/A sky130_fd_sc_hd__or4_4
XFILLER_162_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7465_ _7462_/X _7464_/X _7462_/X _7464_/X vssd1 vssd1 vccd1 vccd1 _7465_/X sky130_fd_sc_hd__a2bb2o_1
X_9204_ _6548_/Y _9809_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9558_/D sky130_fd_sc_hd__mux2_1
X_6416_ _6416_/A vssd1 vssd1 vccd1 vccd1 _6543_/B sky130_fd_sc_hd__inv_2
X_7396_ _7382_/X _7384_/X _7382_/X _7384_/X vssd1 vssd1 vccd1 vccd1 _7396_/X sky130_fd_sc_hd__a2bb2o_1
X_6347_ _6347_/A vssd1 vssd1 vccd1 vccd1 _6347_/Y sky130_fd_sc_hd__inv_2
X_9135_ _9872_/Q _9888_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9135_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9066_ _8041_/Y _8040_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9066_/X sky130_fd_sc_hd__mux2_1
X_6278_ _6275_/X _6277_/Y _6275_/X _6277_/Y vssd1 vssd1 vccd1 vccd1 _6278_/X sky130_fd_sc_hd__o2bb2a_1
X_8017_ _8017_/A _8021_/B vssd1 vssd1 vccd1 vccd1 _8017_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5229_ _9741_/Q vssd1 vssd1 vccd1 vccd1 _5246_/A sky130_fd_sc_hd__inv_2
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9899_ _9903_/CLK _9899_/D vssd1 vssd1 vccd1 vccd1 _9899_/Q sky130_fd_sc_hd__dfxtp_2
X_8919_ _8919_/A _8958_/B _8818_/X vssd1 vssd1 vccd1 vccd1 _8920_/B sky130_fd_sc_hd__or3b_1
XFILLER_169_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5580_ _8177_/A vssd1 vssd1 vccd1 vccd1 _5609_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7250_ _7240_/C _7249_/A _7239_/A _7249_/Y vssd1 vssd1 vccd1 vccd1 _7250_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6201_ _6201_/A vssd1 vssd1 vccd1 vccd1 _6201_/X sky130_fd_sc_hd__buf_1
XFILLER_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7181_ _7171_/C _7180_/A _7170_/A _7180_/Y vssd1 vssd1 vccd1 vccd1 _7181_/X sky130_fd_sc_hd__a22o_1
XFILLER_124_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6132_ _9566_/Q vssd1 vssd1 vccd1 vccd1 _7943_/A sky130_fd_sc_hd__inv_2
XFILLER_85_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6063_ _9858_/Q vssd1 vssd1 vccd1 vccd1 _7986_/A sky130_fd_sc_hd__inv_2
XFILLER_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5014_ _9827_/Q _5011_/X input22/X _5012_/X _5008_/X vssd1 vssd1 vccd1 vccd1 _9827_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9822_ _9929_/CLK _9822_/D vssd1 vssd1 vccd1 vccd1 _9822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9753_ _9796_/CLK _9753_/D vssd1 vssd1 vccd1 vccd1 _9753_/Q sky130_fd_sc_hd__dfxtp_2
X_6965_ _6720_/X _6723_/X _6724_/X _6745_/X vssd1 vssd1 vccd1 vccd1 _6965_/X sky130_fd_sc_hd__o22a_1
XFILLER_81_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8704_ _8703_/A _8703_/B _8703_/X vssd1 vssd1 vccd1 vccd1 _8707_/A sky130_fd_sc_hd__a21bo_1
X_9684_ _9699_/CLK _9684_/D vssd1 vssd1 vccd1 vccd1 _9684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5916_ _5916_/A _9127_/X vssd1 vssd1 vccd1 vccd1 _9595_/D sky130_fd_sc_hd__and2_1
XFILLER_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8635_ _8714_/A _8634_/B _8634_/Y vssd1 vssd1 vccd1 vccd1 _8635_/X sky130_fd_sc_hd__a21o_1
X_6896_ _6896_/A vssd1 vssd1 vccd1 vccd1 _6898_/A sky130_fd_sc_hd__inv_2
XFILLER_179_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5847_ _5847_/A vssd1 vssd1 vccd1 vccd1 _5847_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8566_ _8566_/A _9457_/X vssd1 vssd1 vccd1 vccd1 _8566_/X sky130_fd_sc_hd__or2_1
XFILLER_182_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5778_ _5723_/X _5752_/X _5723_/X _5752_/X vssd1 vssd1 vccd1 vccd1 _5779_/A sky130_fd_sc_hd__a2bb2o_1
X_8497_ _8605_/A _8652_/A _8566_/A _8773_/B vssd1 vssd1 vccd1 vccd1 _8497_/X sky130_fd_sc_hd__o22a_1
XFILLER_147_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7517_ _7210_/A _7137_/Y _7515_/Y _7516_/Y vssd1 vssd1 vccd1 vccd1 _7517_/X sky130_fd_sc_hd__a31o_1
XFILLER_181_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7448_ _7440_/Y _7444_/X _7446_/X _7447_/X vssd1 vssd1 vccd1 vccd1 _7448_/X sky130_fd_sc_hd__o22a_1
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7379_ _7379_/A vssd1 vssd1 vccd1 vccd1 _7398_/B sky130_fd_sc_hd__buf_1
XFILLER_107_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9118_ _9602_/Q _5026_/A _9667_/Q vssd1 vssd1 vccd1 vccd1 _9118_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9049_ _8004_/Y _9048_/X _9052_/S vssd1 vssd1 vccd1 vccd1 _9049_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6750_ _6812_/A _9094_/X _6814_/A _9095_/X vssd1 vssd1 vccd1 vccd1 _6750_/X sky130_fd_sc_hd__or4_4
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5701_ _5701_/A _9635_/Q vssd1 vssd1 vccd1 vccd1 _5704_/B sky130_fd_sc_hd__nor2_2
XFILLER_16_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6681_ _6975_/A _6981_/B _6982_/D _9467_/X vssd1 vssd1 vccd1 vccd1 _6681_/X sky130_fd_sc_hd__or4_4
X_8420_ _9379_/X vssd1 vssd1 vccd1 vccd1 _8580_/B sky130_fd_sc_hd__inv_2
XFILLER_164_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5632_ _5660_/A vssd1 vssd1 vccd1 vccd1 _5632_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8351_ _4790_/X _8333_/Y _8340_/A _8350_/X vssd1 vssd1 vccd1 vccd1 _8351_/X sky130_fd_sc_hd__o22a_1
X_5563_ _5553_/X _5560_/Y _5561_/Y _7651_/A _5557_/X vssd1 vssd1 vccd1 vccd1 _5564_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_191_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7302_ _7302_/A _7302_/B vssd1 vssd1 vccd1 vccd1 _7303_/B sky130_fd_sc_hd__or2_1
X_5494_ _9428_/X _5493_/X _9428_/X _5493_/X vssd1 vssd1 vccd1 vccd1 _5494_/X sky130_fd_sc_hd__a2bb2o_2
X_8282_ _7723_/A _8224_/Y _7738_/A _8222_/X _8281_/X vssd1 vssd1 vccd1 vccd1 _8282_/Y
+ sky130_fd_sc_hd__o221ai_1
X_7233_ _7233_/A _7233_/B vssd1 vssd1 vccd1 vccd1 _7233_/X sky130_fd_sc_hd__or2_1
XFILLER_132_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7164_ _7164_/A _7164_/B vssd1 vssd1 vccd1 vccd1 _7164_/X sky130_fd_sc_hd__or2_1
XFILLER_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6115_ _7083_/B vssd1 vssd1 vccd1 vccd1 _6115_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7095_ _7084_/A _7084_/B _7085_/B vssd1 vssd1 vccd1 vccd1 _7095_/X sky130_fd_sc_hd__a21bo_1
X_6046_ _6018_/Y _6026_/A _6036_/A _6009_/Y _6045_/X vssd1 vssd1 vccd1 vccd1 _6047_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9805_ _9923_/CLK _9805_/D vssd1 vssd1 vccd1 vccd1 _9805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7997_ _7997_/A _8010_/B vssd1 vssd1 vccd1 vccd1 _7997_/Y sky130_fd_sc_hd__nor2_1
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6948_ _5890_/X _6891_/B _6804_/C _6713_/A _6947_/X vssd1 vssd1 vccd1 vccd1 _6948_/X
+ sky130_fd_sc_hd__a41o_1
X_9736_ _9887_/CLK _9736_/D vssd1 vssd1 vccd1 vccd1 _9736_/Q sky130_fd_sc_hd__dfxtp_1
X_6879_ _6865_/X _6867_/X _6865_/X _6867_/X vssd1 vssd1 vccd1 vccd1 _6879_/X sky130_fd_sc_hd__a2bb2o_1
X_9667_ _9858_/CLK _9667_/D vssd1 vssd1 vccd1 vccd1 _9667_/Q sky130_fd_sc_hd__dfxtp_4
X_8618_ _8612_/X _8617_/X _8612_/X _8617_/X vssd1 vssd1 vccd1 vccd1 _8621_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_179_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9598_ _9874_/CLK _9598_/D vssd1 vssd1 vccd1 vccd1 _9598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8549_ _8626_/C _8549_/B vssd1 vssd1 vccd1 vccd1 _8591_/A sky130_fd_sc_hd__nand2_2
XFILLER_194_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _9928_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7920_ _7971_/A _9051_/S _8046_/B vssd1 vssd1 vccd1 vccd1 _7921_/A sky130_fd_sc_hd__or3b_2
X_7851_ _7738_/X _7846_/Y _7673_/B vssd1 vssd1 vccd1 vccd1 _7851_/Y sky130_fd_sc_hd__o21ai_1
X_6802_ _6804_/B vssd1 vssd1 vccd1 vccd1 _6891_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_63_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4994_ _5003_/A vssd1 vssd1 vccd1 vccd1 _4994_/X sky130_fd_sc_hd__clkbuf_2
X_7782_ _8134_/A _7779_/A _7657_/B vssd1 vssd1 vccd1 vccd1 _7782_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_90_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9521_ _9650_/CLK _9521_/D vssd1 vssd1 vccd1 vccd1 _9521_/Q sky130_fd_sc_hd__dfxtp_1
X_6733_ _6723_/C _6732_/A _6722_/A _6732_/Y vssd1 vssd1 vccd1 vccd1 _6733_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6664_ _6659_/X _6663_/X _6659_/X _6663_/X vssd1 vssd1 vccd1 vccd1 _6992_/A sky130_fd_sc_hd__a2bb2o_1
X_9452_ _9451_/X _6353_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _9452_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5615_ _8176_/A _5615_/B vssd1 vssd1 vccd1 vccd1 _9703_/D sky130_fd_sc_hd__nor2_1
X_8403_ _9690_/Q _6561_/Y _8390_/X _8402_/X vssd1 vssd1 vccd1 vccd1 _8403_/X sky130_fd_sc_hd__o22a_1
XFILLER_191_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9383_ _8487_/X _8485_/A _9490_/S vssd1 vssd1 vccd1 vccd1 _9383_/X sky130_fd_sc_hd__mux2_2
X_6595_ _6593_/A _6593_/B _6594_/Y vssd1 vssd1 vccd1 vccd1 _6595_/X sky130_fd_sc_hd__a21o_1
X_8334_ _9551_/Q vssd1 vssd1 vccd1 vccd1 _8334_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5546_ _9420_/X _5469_/X _5554_/A vssd1 vssd1 vccd1 vccd1 _5546_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_151_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8265_ _8123_/A _8249_/X _9903_/Q _8248_/Y _8264_/X vssd1 vssd1 vccd1 vccd1 _8265_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_105_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5477_ _5475_/Y _5476_/Y _5475_/Y _5476_/Y vssd1 vssd1 vccd1 vccd1 _5477_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_132_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7216_ _7522_/A _7283_/B _7490_/A _7238_/B vssd1 vssd1 vccd1 vccd1 _7218_/A sky130_fd_sc_hd__o22a_1
X_8196_ _8211_/B vssd1 vssd1 vccd1 vccd1 _8199_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_132_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7147_ _7147_/A _7147_/B vssd1 vssd1 vccd1 vccd1 _7147_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7078_ _7078_/A _7078_/B vssd1 vssd1 vccd1 vccd1 _7079_/B sky130_fd_sc_hd__or2_1
X_6029_ _6026_/Y _6028_/A _6026_/A _6028_/Y vssd1 vssd1 vccd1 vccd1 _6029_/X sky130_fd_sc_hd__o22a_1
XFILLER_100_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9719_ _9874_/CLK _9719_/D vssd1 vssd1 vccd1 vccd1 _9719_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6380_ _9762_/Q _8229_/A vssd1 vssd1 vccd1 vccd1 _8227_/A sky130_fd_sc_hd__or2_2
X_5400_ _5392_/B _5379_/X _5399_/X _5398_/Y _5364_/A vssd1 vssd1 vccd1 vccd1 _5401_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5331_ _5331_/A _5371_/A vssd1 vssd1 vccd1 vccd1 _5367_/A sky130_fd_sc_hd__or2_1
XFILLER_154_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8050_ _9532_/Q vssd1 vssd1 vccd1 vccd1 _8050_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7001_ _6684_/X _7000_/X _6684_/X _7000_/X vssd1 vssd1 vccd1 vccd1 _7001_/X sky130_fd_sc_hd__a2bb2o_1
X_5262_ _5262_/A vssd1 vssd1 vccd1 vccd1 _9745_/D sky130_fd_sc_hd__inv_2
XFILLER_102_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5193_ _5205_/A vssd1 vssd1 vccd1 vccd1 _5193_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_205_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8952_ _8859_/X _8898_/X _8951_/X vssd1 vssd1 vccd1 vccd1 _8952_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7903_ _7906_/B vssd1 vssd1 vccd1 vccd1 _7903_/Y sky130_fd_sc_hd__inv_2
X_8883_ _8927_/A _8927_/B vssd1 vssd1 vccd1 vccd1 _8883_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7834_ _7713_/X _7829_/Y _7669_/B vssd1 vssd1 vccd1 vccd1 _7834_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_63_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7765_ _9749_/Q vssd1 vssd1 vccd1 vccd1 _7765_/Y sky130_fd_sc_hd__inv_2
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4977_ _4969_/B _9445_/S _4976_/X _4965_/A _4887_/X vssd1 vssd1 vccd1 vccd1 _9845_/D
+ sky130_fd_sc_hd__a221o_1
X_6716_ _6716_/A _6716_/B vssd1 vssd1 vccd1 vccd1 _6716_/X sky130_fd_sc_hd__or2_1
X_9504_ _9503_/X _9635_/Q _9504_/S vssd1 vssd1 vccd1 vccd1 _9504_/X sky130_fd_sc_hd__mux2_1
XPHY_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7696_ _7823_/A vssd1 vssd1 vccd1 vccd1 _7696_/X sky130_fd_sc_hd__buf_2
XFILLER_149_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9435_ _6318_/D _7861_/A _9480_/S vssd1 vssd1 vccd1 vccd1 _9435_/X sky130_fd_sc_hd__mux2_1
X_6647_ _6683_/A _6969_/B _6647_/C vssd1 vssd1 vccd1 vccd1 _6647_/X sky130_fd_sc_hd__or3_4
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6578_ _6578_/A _6578_/B vssd1 vssd1 vccd1 vccd1 _6592_/B sky130_fd_sc_hd__or2_1
X_9366_ _6338_/Y _7726_/X _9480_/S vssd1 vssd1 vccd1 vccd1 _9366_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8317_ _7807_/A _9536_/Q _7803_/A _9535_/Q vssd1 vssd1 vccd1 vccd1 _8369_/D sky130_fd_sc_hd__o22a_1
X_5529_ _5600_/A _5600_/B vssd1 vssd1 vccd1 vccd1 _5599_/A sky130_fd_sc_hd__nand2_1
X_9297_ _9296_/X _7867_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9297_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8248_ _8236_/A _8236_/B _8246_/Y vssd1 vssd1 vccd1 vccd1 _8248_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8179_ _8182_/A _8996_/X vssd1 vssd1 vccd1 vccd1 _9524_/D sky130_fd_sc_hd__or2_1
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _9796_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _9874_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_170_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5880_ _5041_/X _5865_/X _7492_/C _5866_/X _5070_/A vssd1 vssd1 vccd1 vccd1 _9619_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4900_ _5787_/A vssd1 vssd1 vccd1 vccd1 _4900_/X sky130_fd_sc_hd__buf_2
XFILLER_206_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4831_ _9258_/X _4822_/X _7769_/A _4824_/X _4830_/X vssd1 vssd1 vccd1 vccd1 _9905_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4762_ _4834_/A vssd1 vssd1 vccd1 vccd1 _4796_/A sky130_fd_sc_hd__buf_2
X_7550_ _7540_/X _7541_/X _7542_/X _7549_/X vssd1 vssd1 vccd1 vccd1 _7550_/X sky130_fd_sc_hd__o22a_1
X_6501_ _5112_/Y _6427_/A _6492_/X _6499_/Y _6500_/X vssd1 vssd1 vccd1 vccd1 _6501_/Y
+ sky130_fd_sc_hd__o221ai_2
X_7481_ _7428_/X _7480_/X _7428_/X _7480_/X vssd1 vssd1 vccd1 vccd1 _7482_/B sky130_fd_sc_hd__a2bb2o_1
X_9220_ _9825_/Q _7651_/Y _9528_/Q vssd1 vssd1 vccd1 vccd1 _9220_/X sky130_fd_sc_hd__mux2_1
X_6432_ _9795_/Q _6532_/B vssd1 vssd1 vccd1 vccd1 _6432_/Y sky130_fd_sc_hd__nor2_1
X_9151_ _6205_/X input19/X _9155_/S vssd1 vssd1 vccd1 vccd1 _9151_/X sky130_fd_sc_hd__mux2_1
X_6363_ _8184_/A _9751_/Q vssd1 vssd1 vccd1 vccd1 _6363_/Y sky130_fd_sc_hd__nor2_1
X_8102_ _9550_/Q vssd1 vssd1 vccd1 vccd1 _8102_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6294_ _9593_/Q vssd1 vssd1 vccd1 vccd1 _8044_/A sky130_fd_sc_hd__inv_2
XFILLER_114_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9082_ _9081_/X _7850_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9082_/X sky130_fd_sc_hd__mux2_1
X_5314_ _9730_/Q vssd1 vssd1 vccd1 vccd1 _5337_/A sky130_fd_sc_hd__inv_2
X_8033_ _8033_/A _8033_/B vssd1 vssd1 vccd1 vccd1 _8033_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5245_ _5245_/A _5282_/A vssd1 vssd1 vccd1 vccd1 _5278_/A sky130_fd_sc_hd__or2_1
X_5176_ _9769_/Q _5167_/X input29/X _5168_/X _5175_/X vssd1 vssd1 vccd1 vccd1 _9769_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8935_ _8935_/A _9419_/X vssd1 vssd1 vccd1 vccd1 _8935_/X sky130_fd_sc_hd__or2_1
XFILLER_44_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8866_ _8866_/A _8865_/X vssd1 vssd1 vccd1 vccd1 _8866_/X sky130_fd_sc_hd__or2b_1
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8797_ _8797_/A _8797_/B vssd1 vssd1 vccd1 vccd1 _8845_/A sky130_fd_sc_hd__nor2_2
X_7817_ _7755_/X _7812_/Y _7665_/B vssd1 vssd1 vccd1 vccd1 _7817_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_101_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7748_ _8236_/A vssd1 vssd1 vccd1 vccd1 _7748_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7679_ _9922_/Q _7679_/B vssd1 vssd1 vccd1 vccd1 _7879_/A sky130_fd_sc_hd__or2_1
XFILLER_137_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9418_ _9417_/X _6333_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _9418_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9349_ _7621_/X _7585_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9349_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5030_ _5030_/A vssd1 vssd1 vccd1 vccd1 _5030_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6981_ _6981_/A _6981_/B vssd1 vssd1 vccd1 vccd1 _6981_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5932_ _9165_/X _5930_/X _9589_/Q _5931_/X vssd1 vssd1 vccd1 vccd1 _9589_/D sky130_fd_sc_hd__a22o_1
X_8720_ _8875_/A _8800_/B vssd1 vssd1 vccd1 vccd1 _8722_/A sky130_fd_sc_hd__or2_2
XFILLER_179_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8651_ _8650_/A _8650_/B _8699_/A vssd1 vssd1 vccd1 vccd1 _8651_/X sky130_fd_sc_hd__a21bo_1
XFILLER_80_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5863_ _5882_/A _7913_/A vssd1 vssd1 vccd1 vccd1 _5866_/A sky130_fd_sc_hd__or2_2
X_8582_ _8668_/A _8582_/B vssd1 vssd1 vccd1 vccd1 _8589_/A sky130_fd_sc_hd__or2_1
X_5794_ _9674_/Q _9657_/Q _5732_/Y vssd1 vssd1 vccd1 vccd1 _5794_/X sky130_fd_sc_hd__a21o_1
X_4814_ _9911_/Q vssd1 vssd1 vccd1 vccd1 _4814_/X sky130_fd_sc_hd__clkbuf_2
X_7602_ _7602_/A _7602_/B vssd1 vssd1 vccd1 vccd1 _7603_/B sky130_fd_sc_hd__or2_1
XFILLER_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7533_ _7430_/X _7478_/X _7430_/X _7478_/X vssd1 vssd1 vccd1 vccd1 _7533_/X sky130_fd_sc_hd__a2bb2o_1
X_4745_ _4855_/A _4855_/B vssd1 vssd1 vccd1 vccd1 _4929_/C sky130_fd_sc_hd__or2b_1
XFILLER_147_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7464_ _5872_/X _7408_/B _9624_/Q _7321_/D _7463_/X vssd1 vssd1 vccd1 vccd1 _7464_/X
+ sky130_fd_sc_hd__a41o_1
X_9203_ _6547_/Y _9808_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9557_/D sky130_fd_sc_hd__mux2_1
X_6415_ _6413_/Y _6414_/Y _6390_/B vssd1 vssd1 vccd1 vccd1 _6541_/B sky130_fd_sc_hd__o21a_1
X_7395_ _7385_/X _7386_/X _7393_/X _7394_/X vssd1 vssd1 vccd1 vccd1 _7395_/X sky130_fd_sc_hd__o22a_1
X_6346_ _9773_/Q vssd1 vssd1 vccd1 vccd1 _8204_/A sky130_fd_sc_hd__inv_2
XFILLER_134_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9134_ _9871_/Q _9887_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9134_/X sky130_fd_sc_hd__mux2_1
X_9065_ _8039_/X _8038_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9065_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6277_ _6268_/X _6271_/X _6276_/X vssd1 vssd1 vccd1 vccd1 _6277_/Y sky130_fd_sc_hd__o21ai_1
X_8016_ _9002_/X _8022_/B vssd1 vssd1 vccd1 vccd1 _8016_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5228_ _9742_/Q vssd1 vssd1 vccd1 vccd1 _5247_/A sky130_fd_sc_hd__inv_2
X_5159_ _9777_/Q _5155_/X input37/X _5157_/X _5153_/X vssd1 vssd1 vccd1 vccd1 _9777_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9898_ _9898_/CLK _9898_/D vssd1 vssd1 vccd1 vccd1 _9898_/Q sky130_fd_sc_hd__dfxtp_1
X_8918_ _9633_/Q _8916_/Y _5852_/X _8754_/Y _8917_/X vssd1 vssd1 vccd1 vccd1 _8920_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_169_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8849_ _8800_/A _8893_/B _8955_/A _8800_/B vssd1 vssd1 vccd1 vccd1 _8849_/X sky130_fd_sc_hd__o22a_1
XFILLER_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7180_ _7180_/A vssd1 vssd1 vccd1 vccd1 _7180_/Y sky130_fd_sc_hd__inv_2
X_6200_ _6200_/A _6200_/B _6200_/C vssd1 vssd1 vccd1 vccd1 _6203_/A sky130_fd_sc_hd__or3_1
XFILLER_171_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6131_ _6130_/A _6130_/B _6150_/A vssd1 vssd1 vccd1 vccd1 _6131_/X sky130_fd_sc_hd__o21a_1
XFILLER_112_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6062_ _6057_/A _6061_/X _6057_/A _6061_/X vssd1 vssd1 vccd1 vccd1 _6062_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_58_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5013_ _9828_/Q _5011_/X input23/X _5012_/X _5008_/X vssd1 vssd1 vccd1 vccd1 _9828_/D
+ sky130_fd_sc_hd__o221a_1
X_9821_ _9929_/CLK _9821_/D vssd1 vssd1 vccd1 vccd1 _9821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9752_ _9907_/CLK _9752_/D vssd1 vssd1 vccd1 vccd1 _9752_/Q sky130_fd_sc_hd__dfxtp_2
X_6964_ _6964_/A _6964_/B vssd1 vssd1 vccd1 vccd1 _6964_/X sky130_fd_sc_hd__or2_1
XFILLER_81_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8703_ _8703_/A _8703_/B vssd1 vssd1 vccd1 vccd1 _8703_/X sky130_fd_sc_hd__or2_1
X_9683_ _9697_/CLK _9683_/D vssd1 vssd1 vccd1 vccd1 _9683_/Q sky130_fd_sc_hd__dfxtp_4
X_6895_ _6878_/X _6879_/X _6878_/X _6879_/X vssd1 vssd1 vccd1 vccd1 _6896_/A sky130_fd_sc_hd__a2bb2o_1
X_5915_ _5915_/A _9128_/X vssd1 vssd1 vccd1 vccd1 _9596_/D sky130_fd_sc_hd__and2_1
XFILLER_179_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8634_ _8714_/A _8634_/B vssd1 vssd1 vccd1 vccd1 _8634_/Y sky130_fd_sc_hd__nor2_1
X_5846_ _5848_/A vssd1 vssd1 vccd1 vccd1 _5847_/A sky130_fd_sc_hd__inv_2
XFILLER_166_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8565_ _9477_/X vssd1 vssd1 vccd1 vccd1 _8656_/A sky130_fd_sc_hd__inv_2
XFILLER_158_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5777_ _9662_/Q _5774_/X _5769_/X _7110_/A _5772_/X vssd1 vssd1 vccd1 vccd1 _9662_/D
+ sky130_fd_sc_hd__o221a_1
X_8496_ _9381_/X vssd1 vssd1 vccd1 vccd1 _8773_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_182_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7516_ _7210_/A _7137_/Y _7515_/Y vssd1 vssd1 vccd1 vccd1 _7516_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_174_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7447_ _7440_/Y _7444_/X _7440_/Y _7444_/X vssd1 vssd1 vccd1 vccd1 _7447_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_174_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7378_ _7284_/X _7305_/X _7306_/X _7376_/X _7377_/X vssd1 vssd1 vccd1 vccd1 _7378_/X
+ sky130_fd_sc_hd__o221a_1
X_6329_ _6329_/A vssd1 vssd1 vccd1 vccd1 _6486_/B sky130_fd_sc_hd__inv_2
XFILLER_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9117_ _9601_/Q _5029_/A _9667_/Q vssd1 vssd1 vccd1 vccd1 _9117_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9048_ _8005_/Y _9609_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9048_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5700_ _9848_/Q vssd1 vssd1 vccd1 vccd1 _5701_/A sky130_fd_sc_hd__inv_2
XFILLER_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6680_ _6975_/A _6981_/B _6982_/D _9467_/X vssd1 vssd1 vccd1 vccd1 _6682_/A sky130_fd_sc_hd__o22a_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5631_ _5631_/A vssd1 vssd1 vccd1 vccd1 _5631_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8350_ _8340_/C _8349_/X _8345_/X vssd1 vssd1 vccd1 vccd1 _8350_/X sky130_fd_sc_hd__o21a_1
X_5562_ _9713_/Q vssd1 vssd1 vccd1 vccd1 _7651_/A sky130_fd_sc_hd__inv_2
XFILLER_129_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8281_ _7743_/A _8226_/X _7723_/A _8224_/Y _8280_/X vssd1 vssd1 vccd1 vccd1 _8281_/X
+ sky130_fd_sc_hd__a221o_1
X_7301_ _7277_/C _7274_/B _7274_/Y vssd1 vssd1 vccd1 vccd1 _7302_/B sky130_fd_sc_hd__o21ai_1
XFILLER_144_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7232_ _7223_/A _7222_/B _7394_/A _7247_/B _7231_/Y vssd1 vssd1 vccd1 vccd1 _7233_/B
+ sky130_fd_sc_hd__o41a_1
X_5493_ _5491_/Y _5492_/Y _5491_/Y _5492_/Y vssd1 vssd1 vccd1 vccd1 _5493_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7163_ _7195_/A _9430_/X _7156_/A _9431_/X _7162_/Y vssd1 vssd1 vccd1 vccd1 _7164_/B
+ sky130_fd_sc_hd__o41a_1
X_6114_ _6111_/X _6113_/Y _6111_/X _6113_/Y vssd1 vssd1 vccd1 vccd1 _6114_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_86_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7094_ _7085_/A _7085_/B _7086_/B vssd1 vssd1 vccd1 vccd1 _7094_/X sky130_fd_sc_hd__a21bo_1
XFILLER_140_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6045_ _7969_/A _9642_/Q _6034_/Y _6039_/X vssd1 vssd1 vccd1 vccd1 _6045_/X sky130_fd_sc_hd__o22a_2
XFILLER_100_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9804_ _9923_/CLK _9804_/D vssd1 vssd1 vccd1 vccd1 _9804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7996_ _9456_/X _8009_/B vssd1 vssd1 vccd1 vccd1 _7996_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9735_ _9887_/CLK _9735_/D vssd1 vssd1 vccd1 vccd1 _9735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6947_ _6706_/A _6867_/B _6890_/A _6707_/A vssd1 vssd1 vccd1 vccd1 _6947_/X sky130_fd_sc_hd__o22a_1
X_9666_ _9673_/CLK _9666_/D vssd1 vssd1 vccd1 vccd1 _9666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6878_ _6868_/X _6869_/X _6876_/X _6877_/X vssd1 vssd1 vccd1 vccd1 _6878_/X sky130_fd_sc_hd__o22a_1
X_8617_ _8614_/Y _8616_/X _8614_/Y _8616_/X vssd1 vssd1 vccd1 vccd1 _8617_/X sky130_fd_sc_hd__o2bb2a_1
X_5829_ _9644_/Q _5824_/X input47/X _5825_/X _5822_/X vssd1 vssd1 vccd1 vccd1 _9644_/D
+ sky130_fd_sc_hd__o221a_1
X_9597_ _9879_/CLK _9597_/D vssd1 vssd1 vccd1 vccd1 _9597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8548_ _8546_/A _8547_/A _8630_/C _8547_/Y vssd1 vssd1 vccd1 vccd1 _8549_/B sky130_fd_sc_hd__o22a_1
XFILLER_167_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8479_ _8479_/A _8479_/B vssd1 vssd1 vccd1 vccd1 _8479_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7850_ _7723_/X _7848_/B _7839_/X _7849_/Y vssd1 vssd1 vccd1 vccd1 _7850_/Y sky130_fd_sc_hd__a211oi_2
X_6801_ _9427_/X vssd1 vssd1 vccd1 vccd1 _6804_/B sky130_fd_sc_hd__inv_2
XFILLER_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4993_ _9839_/Q _4985_/X input35/X _4987_/X _4991_/X vssd1 vssd1 vccd1 vccd1 _9839_/D
+ sky130_fd_sc_hd__o221a_1
X_7781_ _7781_/A _7781_/B vssd1 vssd1 vccd1 vccd1 _7781_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9520_ _9898_/CLK _9520_/D vssd1 vssd1 vccd1 vccd1 _9521_/D sky130_fd_sc_hd__dfxtp_2
X_6732_ _6732_/A vssd1 vssd1 vccd1 vccd1 _6732_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9451_ _6500_/A _7743_/X _9480_/S vssd1 vssd1 vccd1 vccd1 _9451_/X sky130_fd_sc_hd__mux2_1
X_6663_ _6653_/C _6662_/A _6652_/A _6662_/Y vssd1 vssd1 vccd1 vccd1 _6663_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5614_ _5586_/X _5611_/Y _5612_/Y _7639_/A _5607_/X vssd1 vssd1 vccd1 vccd1 _5615_/B
+ sky130_fd_sc_hd__o32a_1
X_8402_ _8391_/Y _8401_/Y _9689_/Q _8391_/B vssd1 vssd1 vccd1 vccd1 _8402_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_176_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9382_ _8492_/X _8490_/Y _9477_/S vssd1 vssd1 vccd1 vccd1 _9382_/X sky130_fd_sc_hd__mux2_2
X_6594_ _6982_/B vssd1 vssd1 vccd1 vccd1 _6594_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8333_ _9552_/Q vssd1 vssd1 vccd1 vccd1 _8333_/Y sky130_fd_sc_hd__inv_2
X_5545_ _5555_/A _5555_/B vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__nand2_1
XFILLER_144_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8264_ _9902_/Q _8249_/X _8324_/A _8250_/X _8263_/X vssd1 vssd1 vccd1 vccd1 _8264_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_105_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5476_ _5412_/A _5412_/B _5412_/Y vssd1 vssd1 vccd1 vccd1 _5476_/Y sky130_fd_sc_hd__a21oi_1
X_8195_ _8219_/B vssd1 vssd1 vccd1 vccd1 _8211_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_105_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7215_ _9470_/X vssd1 vssd1 vccd1 vccd1 _7238_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_132_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7146_ _7234_/A _7522_/B _7210_/C vssd1 vssd1 vccd1 vccd1 _7147_/B sky130_fd_sc_hd__or3_1
XFILLER_113_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7077_ _7077_/A _7077_/B vssd1 vssd1 vccd1 vccd1 _7078_/B sky130_fd_sc_hd__or2_2
X_6028_ _6028_/A vssd1 vssd1 vccd1 vccd1 _6028_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7979_ _8045_/B vssd1 vssd1 vccd1 vccd1 _8002_/B sky130_fd_sc_hd__buf_2
XFILLER_42_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9718_ _9874_/CLK _9718_/D vssd1 vssd1 vccd1 vccd1 _9718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9649_ _9650_/CLK _9649_/D vssd1 vssd1 vccd1 vccd1 _9649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5330_ _5330_/A _5375_/A vssd1 vssd1 vccd1 vccd1 _5371_/A sky130_fd_sc_hd__or2_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5261_ _5251_/B _5224_/X _5260_/Y _4853_/X _5250_/A vssd1 vssd1 vccd1 vccd1 _5262_/A
+ sky130_fd_sc_hd__o32a_1
X_7000_ _6992_/A _6992_/B _6992_/X vssd1 vssd1 vccd1 vccd1 _7000_/X sky130_fd_sc_hd__a21bo_1
XFILLER_114_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5192_ _5203_/A vssd1 vssd1 vccd1 vccd1 _5192_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8951_ _8892_/X _8893_/X _8894_/Y _8897_/Y vssd1 vssd1 vccd1 vccd1 _8951_/X sky130_fd_sc_hd__o22a_1
X_7902_ _7902_/A _7902_/B vssd1 vssd1 vccd1 vccd1 _7906_/B sky130_fd_sc_hd__or2_1
XFILLER_83_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8882_ _8881_/A _8881_/B _8881_/X vssd1 vssd1 vccd1 vccd1 _8927_/B sky130_fd_sc_hd__a21bo_1
XFILLER_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7833_ _7698_/X _7831_/B _7781_/A _7832_/Y vssd1 vssd1 vccd1 vccd1 _7833_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_63_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7764_ _7761_/X _6335_/A _9914_/Q _6352_/Y _7763_/X vssd1 vssd1 vccd1 vccd1 _7772_/B
+ sky130_fd_sc_hd__o221a_1
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4976_ _9845_/Q vssd1 vssd1 vccd1 vccd1 _4976_/X sky130_fd_sc_hd__buf_2
X_6715_ _6706_/A _6705_/B _6707_/A _6730_/B _6714_/Y vssd1 vssd1 vccd1 vccd1 _6716_/B
+ sky130_fd_sc_hd__o41a_1
X_9503_ _9848_/Q _9667_/Q _9503_/S vssd1 vssd1 vccd1 vccd1 _9503_/X sky130_fd_sc_hd__mux2_1
XPHY_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7695_ _9908_/Q vssd1 vssd1 vccd1 vccd1 _7823_/A sky130_fd_sc_hd__inv_2
XFILLER_192_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _9926_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9434_ _9433_/X _6351_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _9434_/X sky130_fd_sc_hd__mux2_1
X_6646_ _6646_/A _6646_/B vssd1 vssd1 vccd1 vccd1 _6646_/X sky130_fd_sc_hd__or2_1
XFILLER_50_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6577_ _6577_/A _6577_/B vssd1 vssd1 vccd1 vccd1 _6578_/B sky130_fd_sc_hd__or2_1
X_9365_ _7063_/A _7620_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9365_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5528_ _9383_/X _5501_/X _5604_/A vssd1 vssd1 vccd1 vccd1 _5600_/B sky130_fd_sc_hd__o21ai_1
XFILLER_133_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8316_ _4812_/X _8303_/Y _8328_/A _8315_/X vssd1 vssd1 vccd1 vccd1 _8316_/X sky130_fd_sc_hd__o22a_1
XFILLER_3_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9296_ _9769_/Q _9295_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9296_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8247_ _6469_/Y _8246_/Y _8238_/B vssd1 vssd1 vccd1 vccd1 _8247_/X sky130_fd_sc_hd__o21a_1
X_5459_ _9353_/X _9351_/X _5419_/X _5458_/X vssd1 vssd1 vccd1 vccd1 _5483_/A sky130_fd_sc_hd__o22a_1
XFILLER_160_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8178_ _8182_/A _9000_/X vssd1 vssd1 vccd1 vccd1 _9523_/D sky130_fd_sc_hd__or2_1
XFILLER_120_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7129_ _9623_/Q vssd1 vssd1 vccd1 vccd1 _7389_/A sky130_fd_sc_hd__inv_2
XFILLER_115_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4830_ _4830_/A vssd1 vssd1 vccd1 vccd1 _4830_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_159_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4761_ _4836_/A vssd1 vssd1 vccd1 vccd1 _4834_/A sky130_fd_sc_hd__inv_2
X_6500_ _6500_/A _6500_/B vssd1 vssd1 vccd1 vccd1 _6500_/X sky130_fd_sc_hd__or2_1
X_7480_ _7255_/A _7261_/A _7255_/Y vssd1 vssd1 vccd1 vccd1 _7480_/X sky130_fd_sc_hd__a21o_1
XFILLER_146_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6431_ _6429_/Y _6430_/Y _8225_/A vssd1 vssd1 vccd1 vccd1 _6532_/B sky130_fd_sc_hd__o21a_1
X_6362_ _8053_/A vssd1 vssd1 vccd1 vccd1 _8184_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9150_ _6195_/X input18/X _9155_/S vssd1 vssd1 vccd1 vccd1 _9150_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8101_ _9551_/Q _8079_/B _8080_/B vssd1 vssd1 vccd1 vccd1 _8101_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_127_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5313_ _5379_/A vssd1 vssd1 vccd1 vccd1 _5313_/X sky130_fd_sc_hd__clkbuf_2
X_6293_ _6296_/B _6292_/Y _6296_/B _6292_/Y vssd1 vssd1 vccd1 vccd1 _6293_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9081_ _9765_/Q _9080_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9081_/X sky130_fd_sc_hd__mux2_1
X_8032_ _9443_/X _8037_/B vssd1 vssd1 vccd1 vccd1 _8032_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5244_ _5244_/A _5286_/A vssd1 vssd1 vccd1 vccd1 _5282_/A sky130_fd_sc_hd__or2_1
X_5175_ _5660_/A vssd1 vssd1 vccd1 vccd1 _5175_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8934_ _8900_/X _8901_/X _8902_/X _8906_/Y _8865_/X vssd1 vssd1 vccd1 vccd1 _8934_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8865_ _8865_/A _8959_/B _8865_/C vssd1 vssd1 vccd1 vccd1 _8865_/X sky130_fd_sc_hd__or3_1
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7816_ _7726_/X _7814_/B _7781_/A _7815_/Y vssd1 vssd1 vccd1 vccd1 _7816_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8796_ _8796_/A vssd1 vssd1 vccd1 vccd1 _8797_/B sky130_fd_sc_hd__inv_2
XFILLER_24_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7747_ _9922_/Q vssd1 vssd1 vccd1 vccd1 _7882_/A sky130_fd_sc_hd__inv_2
XFILLER_101_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4959_ _9111_/X _4951_/A _9848_/Q _4952_/A _4955_/X vssd1 vssd1 vccd1 vccd1 _9848_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7678_ _9921_/Q _7871_/A vssd1 vssd1 vccd1 vccd1 _7679_/B sky130_fd_sc_hd__or2_1
XFILLER_20_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6629_ _6660_/A _6969_/B _6981_/A _7006_/B vssd1 vssd1 vccd1 vccd1 _6631_/A sky130_fd_sc_hd__o22a_1
X_9417_ _6456_/A _7698_/X _9480_/S vssd1 vssd1 vccd1 vccd1 _9417_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9348_ _7611_/X _7580_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9348_/X sky130_fd_sc_hd__mux2_2
XFILLER_3_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9279_ _7838_/X _9763_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9279_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6980_ _6978_/X _6979_/X _6681_/X _6978_/X vssd1 vssd1 vccd1 vccd1 _6980_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5931_ _5938_/A vssd1 vssd1 vccd1 vccd1 _5931_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8650_ _8650_/A _8650_/B vssd1 vssd1 vccd1 vccd1 _8699_/A sky130_fd_sc_hd__or2_1
X_5862_ _5862_/A _7918_/B vssd1 vssd1 vccd1 vccd1 _7913_/A sky130_fd_sc_hd__or2_4
X_8581_ _8773_/A _8626_/B _7967_/A _8543_/B vssd1 vssd1 vccd1 vccd1 _8582_/B sky130_fd_sc_hd__o22a_1
X_5793_ _8967_/B vssd1 vssd1 vccd1 vccd1 _5793_/X sky130_fd_sc_hd__clkbuf_2
X_4813_ _9282_/X _4809_/X _4812_/X _4810_/X _4806_/X vssd1 vssd1 vccd1 vccd1 _9912_/D
+ sky130_fd_sc_hd__o221a_1
X_7601_ _7601_/A _7601_/B vssd1 vssd1 vccd1 vccd1 _7602_/B sky130_fd_sc_hd__or2_1
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7532_ _7553_/A _7553_/B vssd1 vssd1 vccd1 vccd1 _7532_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4744_ _4744_/A vssd1 vssd1 vccd1 vccd1 _5918_/A sky130_fd_sc_hd__clkinv_4
XFILLER_186_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9202_ _6546_/Y _9807_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9556_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7463_ _7223_/A _7384_/B _7394_/A _7101_/X vssd1 vssd1 vccd1 vccd1 _7463_/X sky130_fd_sc_hd__o22a_1
X_6414_ _8211_/A vssd1 vssd1 vccd1 vccd1 _6414_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7394_ _7394_/A _7400_/B _7394_/C vssd1 vssd1 vccd1 vccd1 _7394_/X sky130_fd_sc_hd__or3_1
X_6345_ _8205_/A vssd1 vssd1 vccd1 vccd1 _6345_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9133_ _9870_/Q _9886_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9133_/X sky130_fd_sc_hd__mux2_1
X_9064_ _8037_/Y _8036_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9064_/X sky130_fd_sc_hd__mux2_1
X_6276_ _8031_/A _6141_/A _8033_/A _6141_/A vssd1 vssd1 vccd1 vccd1 _6276_/X sky130_fd_sc_hd__o22a_1
XFILLER_142_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _9903_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_130_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8015_ _8015_/A _8021_/B vssd1 vssd1 vccd1 vccd1 _8015_/Y sky130_fd_sc_hd__nor2_1
X_5227_ _9743_/Q vssd1 vssd1 vccd1 vccd1 _5248_/A sky130_fd_sc_hd__inv_2
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5158_ _9778_/Q _5155_/X input39/X _5157_/X _5153_/X vssd1 vssd1 vccd1 vccd1 _9778_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5089_ _9802_/Q vssd1 vssd1 vccd1 vccd1 _6318_/B sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_26_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _9656_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8917_ _8958_/A _8955_/B _8959_/A _8821_/B vssd1 vssd1 vccd1 vccd1 _8917_/X sky130_fd_sc_hd__o22a_1
XFILLER_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9897_ _9898_/CLK _9897_/D vssd1 vssd1 vccd1 vccd1 _9897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8848_ _8799_/X _8813_/Y _8814_/X _8815_/X vssd1 vssd1 vccd1 vccd1 _8859_/A sky130_fd_sc_hd__o22a_1
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8779_ _8807_/A _8773_/D _8637_/A _8722_/A _8723_/A vssd1 vssd1 vccd1 vccd1 _8805_/A
+ sky130_fd_sc_hd__o32a_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6130_ _6130_/A _6130_/B vssd1 vssd1 vccd1 vccd1 _6150_/A sky130_fd_sc_hd__nand2_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6061_ _7974_/A _9643_/Q _6048_/A _6045_/X vssd1 vssd1 vccd1 vccd1 _6061_/X sky130_fd_sc_hd__o22a_1
X_5012_ _5030_/A vssd1 vssd1 vccd1 vccd1 _5012_/X sky130_fd_sc_hd__buf_1
XFILLER_38_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9820_ _9929_/CLK _9820_/D vssd1 vssd1 vccd1 vccd1 _9820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9751_ _9819_/CLK _9751_/D vssd1 vssd1 vccd1 vccd1 _9751_/Q sky130_fd_sc_hd__dfxtp_2
X_6963_ _6911_/X _6962_/X _6911_/X _6962_/X vssd1 vssd1 vccd1 vccd1 _6964_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8702_ _8865_/A _8768_/A _8702_/C vssd1 vssd1 vccd1 vccd1 _8703_/B sky130_fd_sc_hd__or3_1
XFILLER_179_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9682_ _9697_/CLK _9682_/D vssd1 vssd1 vccd1 vccd1 _9682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5914_ _5915_/A _9129_/X vssd1 vssd1 vccd1 vccd1 _9597_/D sky130_fd_sc_hd__and2_1
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6894_ _6889_/X _6893_/X _6889_/X _6893_/X vssd1 vssd1 vccd1 vccd1 _6926_/A sky130_fd_sc_hd__a2bb2o_1
X_8633_ _8633_/A _8715_/A vssd1 vssd1 vccd1 vccd1 _8634_/B sky130_fd_sc_hd__nor2_2
X_5845_ _5882_/A _7912_/A vssd1 vssd1 vccd1 vccd1 _5848_/A sky130_fd_sc_hd__or2_4
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8564_ _8564_/A _8563_/X vssd1 vssd1 vccd1 vccd1 _8571_/A sky130_fd_sc_hd__or2b_1
X_5776_ _5776_/A vssd1 vssd1 vccd1 vccd1 _7110_/A sky130_fd_sc_hd__inv_2
X_8495_ _8495_/A vssd1 vssd1 vccd1 vccd1 _8536_/C sky130_fd_sc_hd__inv_2
X_7515_ _7498_/X _7508_/X _7509_/X _7514_/X vssd1 vssd1 vccd1 vccd1 _7515_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_107_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7446_ _5872_/X _7291_/B _7210_/A _7359_/Y _7445_/X vssd1 vssd1 vccd1 vccd1 _7446_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_162_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7377_ _7264_/X _7265_/X _7280_/X _7283_/X vssd1 vssd1 vccd1 vccd1 _7377_/X sky130_fd_sc_hd__o22a_1
X_9116_ _9600_/Q _5032_/A _9667_/Q vssd1 vssd1 vccd1 vccd1 _9116_/X sky130_fd_sc_hd__mux2_1
X_6328_ _8056_/A _5218_/X _6327_/Y vssd1 vssd1 vccd1 vccd1 _6329_/A sky130_fd_sc_hd__a21oi_2
XFILLER_143_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6259_ _9586_/Q vssd1 vssd1 vccd1 vccd1 _8029_/A sky130_fd_sc_hd__inv_2
XFILLER_107_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9047_ _8002_/Y _9046_/X _9053_/S vssd1 vssd1 vccd1 vccd1 _9047_/X sky130_fd_sc_hd__mux2_2
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5630_ _8176_/A _5630_/B vssd1 vssd1 vccd1 vccd1 _9700_/D sky130_fd_sc_hd__nor2_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5561_ _5561_/A _5561_/B vssd1 vssd1 vccd1 vccd1 _5561_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8280_ _7743_/A _8226_/X _8279_/X vssd1 vssd1 vccd1 vccd1 _8280_/X sky130_fd_sc_hd__o21a_1
X_7300_ _7288_/A _7288_/B _7372_/A vssd1 vssd1 vccd1 vccd1 _7303_/A sky130_fd_sc_hd__a21o_1
X_5492_ _5423_/A _5423_/B _5423_/Y vssd1 vssd1 vccd1 vccd1 _5492_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_156_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7231_ _7234_/C _7231_/B vssd1 vssd1 vccd1 vccd1 _7231_/Y sky130_fd_sc_hd__nand2_1
XFILLER_144_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7162_ _7165_/C _7162_/B vssd1 vssd1 vccd1 vccd1 _7162_/Y sky130_fd_sc_hd__nand2_1
XFILLER_140_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6113_ _8003_/A _9649_/Q _6103_/X _6104_/X vssd1 vssd1 vccd1 vccd1 _6113_/Y sky130_fd_sc_hd__o22ai_1
X_7093_ _7086_/A _7086_/B _7087_/B vssd1 vssd1 vccd1 vccd1 _7093_/X sky130_fd_sc_hd__a21bo_1
XFILLER_140_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6044_ _9855_/Q vssd1 vssd1 vccd1 vccd1 _7969_/A sky130_fd_sc_hd__inv_2
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9803_ _9923_/CLK _9803_/D vssd1 vssd1 vccd1 vccd1 _9803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7995_ _7995_/A _8003_/B vssd1 vssd1 vccd1 vccd1 _7995_/X sky130_fd_sc_hd__or2_1
XFILLER_81_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9734_ _9893_/CLK _9734_/D vssd1 vssd1 vccd1 vccd1 _9734_/Q sky130_fd_sc_hd__dfxtp_1
X_6946_ _6849_/X _6851_/X _6849_/X _6851_/X vssd1 vssd1 vccd1 vccd1 _6946_/X sky130_fd_sc_hd__a2bb2o_1
X_9665_ _9715_/CLK _9665_/D vssd1 vssd1 vccd1 vccd1 _9665_/Q sky130_fd_sc_hd__dfxtp_1
X_6877_ _6877_/A _6883_/B _6877_/C vssd1 vssd1 vccd1 vccd1 _6877_/X sky130_fd_sc_hd__or3_1
X_8616_ _8735_/A _8768_/A _8535_/X vssd1 vssd1 vccd1 vccd1 _8616_/X sky130_fd_sc_hd__or3b_1
XFILLER_194_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5828_ _9645_/Q _5824_/X input17/X _5825_/X _5822_/X vssd1 vssd1 vccd1 vccd1 _9645_/D
+ sky130_fd_sc_hd__o221a_1
X_9596_ _9879_/CLK _9596_/D vssd1 vssd1 vccd1 vccd1 _9596_/Q sky130_fd_sc_hd__dfxtp_1
X_8547_ _8547_/A vssd1 vssd1 vccd1 vccd1 _8547_/Y sky130_fd_sc_hd__inv_2
X_5759_ _6982_/C _9666_/Q _6982_/C _9666_/Q vssd1 vssd1 vccd1 vccd1 _5759_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_194_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8478_ _8478_/A _8531_/A vssd1 vssd1 vccd1 vccd1 _8479_/B sky130_fd_sc_hd__nor2_2
XFILLER_135_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7429_ _7428_/A _7428_/B _7428_/X vssd1 vssd1 vccd1 vccd1 _7429_/X sky130_fd_sc_hd__a21bo_1
XFILLER_78_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6800_ _6800_/A _6862_/A vssd1 vssd1 vccd1 vccd1 _6807_/C sky130_fd_sc_hd__nor2_2
X_4992_ _9840_/Q _4985_/X input36/X _4987_/X _4991_/X vssd1 vssd1 vccd1 vccd1 _9840_/D
+ sky130_fd_sc_hd__o221a_1
X_7780_ _7780_/A vssd1 vssd1 vccd1 vccd1 _7781_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_90_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6731_ _9618_/Q _6774_/B _6742_/A vssd1 vssd1 vccd1 vccd1 _6732_/A sky130_fd_sc_hd__and3_1
X_6662_ _6662_/A vssd1 vssd1 vccd1 vccd1 _6662_/Y sky130_fd_sc_hd__inv_2
X_9450_ _9449_/X _6335_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _9450_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5613_ _9703_/Q vssd1 vssd1 vccd1 vccd1 _7639_/A sky130_fd_sc_hd__inv_2
X_9381_ _8468_/X _8466_/A _9477_/S vssd1 vssd1 vccd1 vccd1 _9381_/X sky130_fd_sc_hd__mux2_2
X_8401_ _9688_/Q _6564_/X _8392_/X _8400_/X vssd1 vssd1 vccd1 vccd1 _8401_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_31_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8332_ _7807_/A _9536_/Q _8369_/D _8327_/X _8375_/B vssd1 vssd1 vccd1 vccd1 _8332_/Y
+ sky130_fd_sc_hd__a221oi_2
X_6593_ _6593_/A _6593_/B vssd1 vssd1 vccd1 vccd1 _6982_/B sky130_fd_sc_hd__or2_2
XFILLER_191_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5544_ _9421_/X _5473_/X _5560_/A vssd1 vssd1 vccd1 vccd1 _5555_/B sky130_fd_sc_hd__o21ai_1
X_8263_ _7657_/A _8259_/Y _9901_/Q _8250_/X _8262_/Y vssd1 vssd1 vccd1 vccd1 _8263_/X
+ sky130_fd_sc_hd__o221a_1
X_5475_ _5475_/A vssd1 vssd1 vccd1 vccd1 _5475_/Y sky130_fd_sc_hd__inv_2
X_8194_ _8227_/B vssd1 vssd1 vccd1 vccd1 _8219_/B sky130_fd_sc_hd__clkbuf_2
X_7214_ _7400_/A vssd1 vssd1 vccd1 vccd1 _7490_/A sky130_fd_sc_hd__buf_4
X_7145_ _7145_/A vssd1 vssd1 vccd1 vccd1 _7210_/C sky130_fd_sc_hd__inv_2
XFILLER_113_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7076_ _7076_/A _7076_/B vssd1 vssd1 vccd1 vccd1 _7077_/B sky130_fd_sc_hd__or2_1
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6027_ _9853_/Q _6014_/B _6019_/Y _6017_/B vssd1 vssd1 vccd1 vccd1 _6028_/A sky130_fd_sc_hd__o22a_1
XFILLER_39_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7978_ _8025_/A vssd1 vssd1 vccd1 vccd1 _8045_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_42_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _5890_/X _6774_/B _6713_/A _6842_/Y _6928_/X vssd1 vssd1 vccd1 vccd1 _6929_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_81_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9717_ _9874_/CLK _9717_/D vssd1 vssd1 vccd1 vccd1 _9717_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9648_ _9828_/CLK _9648_/D vssd1 vssd1 vccd1 vccd1 _9648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9579_ _9910_/CLK _9579_/D vssd1 vssd1 vccd1 vccd1 _9579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5260_ _9745_/Q _5260_/B vssd1 vssd1 vccd1 vccd1 _5260_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5191_ _6331_/A _5203_/A input21/X _5205_/A _5187_/X vssd1 vssd1 vccd1 vccd1 _9762_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_141_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8950_ _8899_/X _8925_/X _8926_/X _8928_/Y vssd1 vssd1 vccd1 vccd1 _8950_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_110_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7901_ _7901_/A vssd1 vssd1 vccd1 vccd1 _7902_/A sky130_fd_sc_hd__buf_2
XFILLER_209_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8881_ _8881_/A _8881_/B vssd1 vssd1 vccd1 vccd1 _8881_/X sky130_fd_sc_hd__or2_1
X_7832_ _7835_/B vssd1 vssd1 vccd1 vccd1 _7832_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7763_ _7778_/B _9748_/Q _7869_/A _9770_/Q vssd1 vssd1 vccd1 vccd1 _7763_/X sky130_fd_sc_hd__o22a_2
X_4975_ _4965_/A _4972_/Y _4973_/X _9445_/S _4974_/X vssd1 vssd1 vccd1 vccd1 _9846_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_189_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6714_ _6717_/C _6714_/B vssd1 vssd1 vccd1 vccd1 _6714_/Y sky130_fd_sc_hd__nand2_1
X_9502_ _9501_/X _7006_/A _9507_/S vssd1 vssd1 vccd1 vccd1 _9502_/X sky130_fd_sc_hd__mux2_1
XPHY_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7694_ _4790_/X _6413_/Y _8324_/A _8191_/A _7693_/X vssd1 vssd1 vccd1 vccd1 _7705_/B
+ sky130_fd_sc_hd__o221a_1
X_9433_ _5108_/Y _7738_/X _9480_/S vssd1 vssd1 vccd1 vccd1 _9433_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6645_ _6678_/A _9463_/X _6683_/A _9464_/X _6644_/Y vssd1 vssd1 vccd1 vccd1 _6646_/B
+ sky130_fd_sc_hd__o41a_1
X_6576_ _6576_/A _6576_/B vssd1 vssd1 vccd1 vccd1 _6577_/B sky130_fd_sc_hd__or2_1
X_9364_ _7625_/X _7587_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9364_/X sky130_fd_sc_hd__mux2_1
X_5527_ _5605_/A _5605_/B vssd1 vssd1 vccd1 vccd1 _5604_/A sky130_fd_sc_hd__nand2_1
X_9295_ _7864_/X _9769_/Q _9327_/S vssd1 vssd1 vccd1 vccd1 _9295_/X sky130_fd_sc_hd__mux2_1
X_8315_ _8328_/C _8313_/X _8314_/X vssd1 vssd1 vccd1 vccd1 _8315_/X sky130_fd_sc_hd__o21a_1
X_8246_ _8246_/A vssd1 vssd1 vccd1 vccd1 _8246_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5458_ _9359_/X _9358_/X _5420_/X _5457_/X vssd1 vssd1 vccd1 vccd1 _5458_/X sky130_fd_sc_hd__o22a_1
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8177_ _8177_/A vssd1 vssd1 vccd1 vccd1 _8182_/A sky130_fd_sc_hd__buf_1
X_5389_ _9720_/Q _5389_/B vssd1 vssd1 vccd1 vccd1 _5389_/Y sky130_fd_sc_hd__nor2_1
X_7128_ _7247_/A vssd1 vssd1 vccd1 vccd1 _7522_/A sky130_fd_sc_hd__buf_2
XFILLER_59_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7059_ _7059_/A vssd1 vssd1 vccd1 vccd1 _7078_/A sky130_fd_sc_hd__inv_2
XFILLER_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4760_ _9525_/D _9282_/S vssd1 vssd1 vccd1 vccd1 _4836_/A sky130_fd_sc_hd__or2_4
XFILLER_174_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6430_ _8227_/A vssd1 vssd1 vccd1 vccd1 _6430_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6361_ _9846_/Q vssd1 vssd1 vccd1 vccd1 _8053_/A sky130_fd_sc_hd__inv_2
X_8100_ _9552_/Q _8080_/B _8081_/B vssd1 vssd1 vccd1 vccd1 _8100_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_115_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5312_ _9335_/X _5348_/B vssd1 vssd1 vccd1 vccd1 _5379_/A sky130_fd_sc_hd__or2_1
X_6292_ _8040_/A _6193_/X _6296_/A vssd1 vssd1 vccd1 vccd1 _6292_/Y sky130_fd_sc_hd__o21ai_1
X_9080_ _7847_/X _9765_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9080_/X sky130_fd_sc_hd__mux2_1
X_8031_ _8031_/A _8033_/B vssd1 vssd1 vccd1 vccd1 _8031_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5243_ _5243_/A _5290_/A vssd1 vssd1 vccd1 vccd1 _5286_/A sky130_fd_sc_hd__or2_1
X_5174_ _5790_/A vssd1 vssd1 vccd1 vccd1 _5660_/A sky130_fd_sc_hd__buf_2
XFILLER_102_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8933_ _8919_/A _8821_/B _8878_/A _8754_/Y _8876_/A vssd1 vssd1 vccd1 vccd1 _8933_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_83_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8864_ _8938_/A _9396_/X _8865_/A _8821_/B vssd1 vssd1 vccd1 vccd1 _8866_/A sky130_fd_sc_hd__o22a_1
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7815_ _7819_/B vssd1 vssd1 vccd1 vccd1 _7815_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8795_ _8382_/X _8408_/X _8382_/X _8408_/X vssd1 vssd1 vccd1 vccd1 _8796_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_200_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7746_ _4786_/X _8204_/A _9913_/Q _6353_/Y _7745_/X vssd1 vssd1 vccd1 vccd1 _7752_/C
+ sky130_fd_sc_hd__o221a_1
X_4958_ _9112_/X _4951_/X _9849_/Q _4952_/X _4955_/X vssd1 vssd1 vccd1 vccd1 _9849_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7677_ _9920_/Q _7677_/B vssd1 vssd1 vccd1 vccd1 _7871_/A sky130_fd_sc_hd__or2_1
X_4889_ _9734_/Q _4865_/X _9882_/Q _4866_/X _4887_/X vssd1 vssd1 vccd1 vccd1 _9882_/D
+ sky130_fd_sc_hd__a221o_1
X_9416_ _8523_/X _8521_/A _9490_/S vssd1 vssd1 vccd1 vccd1 _9416_/X sky130_fd_sc_hd__mux2_2
X_6628_ _6766_/A vssd1 vssd1 vccd1 vccd1 _6981_/A sky130_fd_sc_hd__buf_2
XFILLER_20_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9347_ _7631_/Y _7592_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9347_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6559_ _6575_/B vssd1 vssd1 vccd1 vccd1 _6559_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9278_ _9277_/X input21/X _9282_/S vssd1 vssd1 vccd1 vccd1 _9278_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8229_ _8229_/A _8231_/B vssd1 vssd1 vccd1 vccd1 _8229_/X sky130_fd_sc_hd__or2_1
XFILLER_160_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_7_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _9924_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_93_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5930_ _5937_/A vssd1 vssd1 vccd1 vccd1 _5930_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5861_ _5860_/X _5847_/A _5041_/A _5848_/A _5853_/X vssd1 vssd1 vccd1 vccd1 _9627_/D
+ sky130_fd_sc_hd__o221a_1
X_7600_ _7600_/A _7600_/B vssd1 vssd1 vccd1 vccd1 _7601_/B sky130_fd_sc_hd__or2_1
XFILLER_194_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8580_ _9634_/Q _8580_/B _8626_/C vssd1 vssd1 vccd1 vccd1 _8668_/A sky130_fd_sc_hd__and3_1
X_5792_ _9658_/Q _5774_/X _5787_/X _7089_/A _5791_/X vssd1 vssd1 vccd1 vccd1 _9658_/D
+ sky130_fd_sc_hd__o221a_1
X_4812_ _9912_/Q vssd1 vssd1 vccd1 vccd1 _4812_/X sky130_fd_sc_hd__buf_2
XFILLER_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4743_ _5128_/A vssd1 vssd1 vccd1 vccd1 _4743_/X sky130_fd_sc_hd__clkbuf_2
X_7531_ _7514_/A _7514_/B _7514_/X vssd1 vssd1 vccd1 vccd1 _7553_/B sky130_fd_sc_hd__a21bo_1
X_7462_ _7367_/X _7368_/X _7367_/X _7368_/X vssd1 vssd1 vccd1 vccd1 _7462_/X sky130_fd_sc_hd__a2bb2o_1
X_9201_ _6545_/Y _9806_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9555_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6413_ _9771_/Q vssd1 vssd1 vccd1 vccd1 _6413_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7393_ _7393_/A _7393_/B vssd1 vssd1 vccd1 vccd1 _7393_/X sky130_fd_sc_hd__or2_1
X_6344_ _9776_/Q vssd1 vssd1 vccd1 vccd1 _6344_/Y sky130_fd_sc_hd__inv_2
X_9132_ _9869_/Q _9885_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9132_/X sky130_fd_sc_hd__mux2_1
X_6275_ _8036_/A _6140_/A _9589_/Q _6170_/A vssd1 vssd1 vccd1 vccd1 _6275_/X sky130_fd_sc_hd__o22a_1
X_9063_ _8034_/Y _8033_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9063_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8014_ _9452_/X _8022_/B vssd1 vssd1 vccd1 vccd1 _8014_/Y sky130_fd_sc_hd__nor2_1
X_5226_ _9744_/Q vssd1 vssd1 vccd1 vccd1 _5249_/A sky130_fd_sc_hd__inv_2
X_5157_ _5205_/A vssd1 vssd1 vccd1 vccd1 _5157_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5088_ _5092_/A _5088_/B vssd1 vssd1 vccd1 vccd1 _9803_/D sky130_fd_sc_hd__nor2_1
XFILLER_56_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8916_ _8955_/B vssd1 vssd1 vccd1 vccd1 _8916_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9896_ _9930_/CLK _9896_/D vssd1 vssd1 vccd1 vccd1 _9896_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8847_ _8816_/X _8836_/X _8837_/X _8838_/X vssd1 vssd1 vccd1 vccd1 _8847_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8778_ _5852_/X _8656_/X _8776_/X _8777_/Y vssd1 vssd1 vccd1 vccd1 _8778_/X sky130_fd_sc_hd__a31o_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7729_ _7728_/X _9771_/Q _7692_/X _5181_/X vssd1 vssd1 vccd1 vccd1 _7729_/X sky130_fd_sc_hd__o22a_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6060_ _6057_/Y _6059_/A _6057_/A _6059_/Y vssd1 vssd1 vccd1 vccd1 _6060_/X sky130_fd_sc_hd__o22a_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5011_ _5028_/A vssd1 vssd1 vccd1 vccd1 _5011_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9750_ _9750_/CLK _9750_/D vssd1 vssd1 vccd1 vccd1 _9750_/Q sky130_fd_sc_hd__dfxtp_1
X_6962_ _6738_/A _6744_/A _6738_/Y vssd1 vssd1 vccd1 vccd1 _6962_/X sky130_fd_sc_hd__a21o_1
XFILLER_93_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8701_ _8563_/X _8659_/X _8660_/X _8661_/X vssd1 vssd1 vccd1 vccd1 _8703_/A sky130_fd_sc_hd__o22a_1
XFILLER_179_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9681_ _9699_/CLK _9681_/D vssd1 vssd1 vccd1 vccd1 _9681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5913_ _5915_/A _9130_/X vssd1 vssd1 vccd1 vccd1 _9598_/D sky130_fd_sc_hd__and2_1
X_6893_ _6883_/C _6892_/A _6882_/A _6892_/Y vssd1 vssd1 vccd1 vccd1 _6893_/X sky130_fd_sc_hd__a22o_1
X_8632_ _8627_/X _8631_/X _8627_/X _8631_/X vssd1 vssd1 vccd1 vccd1 _8714_/A sky130_fd_sc_hd__a2bb2o_2
X_5844_ _5844_/A _5862_/A vssd1 vssd1 vccd1 vccd1 _7912_/A sky130_fd_sc_hd__or2_4
X_8563_ _8576_/A _8652_/A _8610_/C vssd1 vssd1 vccd1 vccd1 _8563_/X sky130_fd_sc_hd__or3_4
XFILLER_21_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5775_ _5719_/X _5753_/X _5719_/X _5753_/X vssd1 vssd1 vccd1 vccd1 _5776_/A sky130_fd_sc_hd__a2bb2o_1
X_7514_ _7514_/A _7514_/B vssd1 vssd1 vccd1 vccd1 _7514_/X sky130_fd_sc_hd__or2_2
XFILLER_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8494_ _8652_/A vssd1 vssd1 vccd1 vccd1 _8610_/B sky130_fd_sc_hd__inv_2
XFILLER_159_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7445_ _7494_/A _7222_/B _7234_/A _7247_/B vssd1 vssd1 vccd1 vccd1 _7445_/X sky130_fd_sc_hd__o22a_1
XFILLER_107_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7376_ _7376_/A _7376_/B vssd1 vssd1 vccd1 vccd1 _7376_/X sky130_fd_sc_hd__or2_1
X_6327_ _8056_/A _9749_/Q vssd1 vssd1 vccd1 vccd1 _6327_/Y sky130_fd_sc_hd__nor2_2
X_9115_ _9599_/Q _4978_/A _9667_/Q vssd1 vssd1 vccd1 vccd1 _9115_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6258_ _6265_/C _6257_/X _6265_/C _6257_/X vssd1 vssd1 vccd1 vccd1 _6258_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9046_ _8000_/Y _9045_/X _9052_/S vssd1 vssd1 vccd1 vccd1 _9046_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5209_ _9754_/Q vssd1 vssd1 vccd1 vccd1 _8236_/A sky130_fd_sc_hd__buf_2
XFILLER_69_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6189_ _6200_/C _6189_/B vssd1 vssd1 vccd1 vccd1 _6189_/X sky130_fd_sc_hd__and2_1
XFILLER_123_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9879_ _9879_/CLK _9879_/D vssd1 vssd1 vccd1 vccd1 _9879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_10_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _9898_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5560_ _5560_/A vssd1 vssd1 vccd1 vccd1 _5560_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5491_ _5491_/A vssd1 vssd1 vccd1 vccd1 _5491_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _9673_/CLK sky130_fd_sc_hd__clkbuf_16
X_7230_ _9624_/Q _7291_/B _7230_/C vssd1 vssd1 vccd1 vccd1 _7231_/B sky130_fd_sc_hd__and3_1
XFILLER_171_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7161_ _7273_/A _7210_/B _7548_/A vssd1 vssd1 vccd1 vccd1 _7162_/B sky130_fd_sc_hd__and3_1
X_6112_ _6108_/X _6111_/X _6108_/X _6111_/X vssd1 vssd1 vccd1 vccd1 _6112_/X sky130_fd_sc_hd__o2bb2a_1
X_7092_ _7087_/A _7087_/B _7088_/B vssd1 vssd1 vccd1 vccd1 _7092_/X sky130_fd_sc_hd__a21bo_1
XFILLER_140_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6043_ _9856_/Q _6041_/Y _7974_/A _9643_/Q vssd1 vssd1 vccd1 vccd1 _6048_/A sky130_fd_sc_hd__a22o_1
XFILLER_100_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9802_ _9923_/CLK _9802_/D vssd1 vssd1 vccd1 vccd1 _9802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7994_ _8992_/X _8030_/B vssd1 vssd1 vccd1 vccd1 _7994_/X sky130_fd_sc_hd__and2_1
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9733_ _9895_/CLK _9733_/D vssd1 vssd1 vccd1 vccd1 _9733_/Q sky130_fd_sc_hd__dfxtp_1
X_6945_ _6943_/X _6944_/X _6943_/X _6944_/X vssd1 vssd1 vccd1 vccd1 _6945_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_179_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9664_ _9673_/CLK _9664_/D vssd1 vssd1 vccd1 vccd1 _9664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6876_ _6876_/A _6876_/B vssd1 vssd1 vccd1 vccd1 _6876_/X sky130_fd_sc_hd__or2_1
XFILLER_194_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8615_ _9477_/X vssd1 vssd1 vccd1 vccd1 _8768_/A sky130_fd_sc_hd__clkbuf_2
X_5827_ _9646_/Q _5824_/X input18/X _5825_/X _5822_/X vssd1 vssd1 vccd1 vccd1 _9646_/D
+ sky130_fd_sc_hd__o221a_1
X_9595_ _9930_/CLK _9595_/D vssd1 vssd1 vccd1 vccd1 _9595_/Q sky130_fd_sc_hd__dfxtp_1
X_8546_ _8546_/A vssd1 vssd1 vccd1 vccd1 _8630_/C sky130_fd_sc_hd__inv_2
X_5758_ _9683_/Q vssd1 vssd1 vccd1 vccd1 _6982_/C sky130_fd_sc_hd__inv_2
X_8477_ _8473_/X _8476_/X _8473_/X _8476_/X vssd1 vssd1 vccd1 vccd1 _8479_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_163_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5689_ _5689_/A vssd1 vssd1 vccd1 vccd1 _5689_/X sky130_fd_sc_hd__clkbuf_2
X_7428_ _7428_/A _7428_/B vssd1 vssd1 vccd1 vccd1 _7428_/X sky130_fd_sc_hd__or2_1
XFILLER_190_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7359_ _7359_/A vssd1 vssd1 vccd1 vccd1 _7359_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9029_ _7973_/Y _9602_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9029_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4991_ _4991_/A vssd1 vssd1 vccd1 vccd1 _4991_/X sky130_fd_sc_hd__buf_2
XFILLER_90_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6730_ _6730_/A _6730_/B vssd1 vssd1 vccd1 vccd1 _6742_/A sky130_fd_sc_hd__or2_1
XFILLER_149_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6661_ _9614_/Q _6691_/B _6672_/A vssd1 vssd1 vccd1 vccd1 _6662_/A sky130_fd_sc_hd__and3_1
X_9380_ _8464_/X _8462_/Y _9490_/S vssd1 vssd1 vccd1 vccd1 _9380_/X sky130_fd_sc_hd__mux2_2
X_5612_ _5612_/A _5612_/B vssd1 vssd1 vccd1 vccd1 _5612_/Y sky130_fd_sc_hd__nor2_1
X_6592_ _6596_/A _6592_/B vssd1 vssd1 vccd1 vccd1 _6593_/B sky130_fd_sc_hd__or2_1
X_8400_ _9687_/Q _6567_/Y _8394_/Y _8399_/X vssd1 vssd1 vccd1 vccd1 _8400_/X sky130_fd_sc_hd__o22a_1
X_5543_ _5561_/A _5561_/B vssd1 vssd1 vccd1 vccd1 _5560_/A sky130_fd_sc_hd__nand2_1
X_8331_ _8331_/A _8331_/B _8330_/X _8314_/X vssd1 vssd1 vccd1 vccd1 _8375_/B sky130_fd_sc_hd__or4bb_4
XFILLER_191_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8262_ _7788_/A _8259_/A _8261_/X vssd1 vssd1 vccd1 vccd1 _8262_/Y sky130_fd_sc_hd__o21ai_1
X_5474_ _9421_/X _5473_/X _9421_/X _5473_/X vssd1 vssd1 vccd1 vccd1 _5561_/A sky130_fd_sc_hd__a2bb2oi_1
XFILLER_117_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8193_ _8231_/B vssd1 vssd1 vccd1 vccd1 _8227_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_117_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7213_ _7384_/C vssd1 vssd1 vccd1 vccd1 _7400_/A sky130_fd_sc_hd__clkbuf_2
X_7144_ _7223_/A _7178_/B vssd1 vssd1 vccd1 vccd1 _7145_/A sky130_fd_sc_hd__or2_2
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7075_ _7075_/A _7075_/B vssd1 vssd1 vccd1 vccd1 _7076_/B sky130_fd_sc_hd__or2_1
X_6026_ _6026_/A vssd1 vssd1 vccd1 vccd1 _6026_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7977_ _8047_/B vssd1 vssd1 vccd1 vccd1 _8025_/A sky130_fd_sc_hd__inv_2
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6928_ _6706_/A _6705_/B _6707_/A _6730_/B vssd1 vssd1 vccd1 vccd1 _6928_/X sky130_fd_sc_hd__o22a_1
X_9716_ _9874_/CLK _9716_/D vssd1 vssd1 vccd1 vccd1 _9716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9647_ _9650_/CLK _9647_/D vssd1 vssd1 vccd1 vccd1 _9647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6859_ _6859_/A _6859_/B vssd1 vssd1 vccd1 vccd1 _6859_/X sky130_fd_sc_hd__or2_2
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9578_ _9578_/CLK _9578_/D vssd1 vssd1 vccd1 vccd1 _9578_/Q sky130_fd_sc_hd__dfxtp_1
X_8529_ _8576_/A _8584_/B _8529_/C vssd1 vssd1 vccd1 vccd1 _8529_/X sky130_fd_sc_hd__or3_1
XFILLER_148_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5190_ _9762_/Q vssd1 vssd1 vccd1 vccd1 _6331_/A sky130_fd_sc_hd__buf_2
XFILLER_205_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7900_ _7683_/A _7683_/B _7899_/Y vssd1 vssd1 vccd1 vccd1 _7900_/X sky130_fd_sc_hd__a21o_1
X_8880_ _8820_/X _8834_/X _8818_/X _8835_/X vssd1 vssd1 vccd1 vccd1 _8881_/B sky130_fd_sc_hd__o22a_1
XFILLER_36_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7831_ _7831_/A _7831_/B vssd1 vssd1 vccd1 vccd1 _7835_/B sky130_fd_sc_hd__or2_1
X_4974_ _4991_/A vssd1 vssd1 vccd1 vccd1 _4974_/X sky130_fd_sc_hd__clkbuf_4
X_7762_ _9919_/Q vssd1 vssd1 vccd1 vccd1 _7869_/A sky130_fd_sc_hd__inv_2
XFILLER_24_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7693_ _7692_/X _5181_/X _9907_/Q _6337_/Y vssd1 vssd1 vccd1 vccd1 _7693_/X sky130_fd_sc_hd__o2bb2a_1
X_9501_ _9500_/X _7234_/A _9506_/S vssd1 vssd1 vccd1 vccd1 _9501_/X sky130_fd_sc_hd__mux2_1
X_6713_ _6713_/A _6774_/B _6713_/C vssd1 vssd1 vccd1 vccd1 _6714_/B sky130_fd_sc_hd__and3_1
XFILLER_177_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6644_ _6647_/C _6644_/B vssd1 vssd1 vccd1 vccd1 _6644_/Y sky130_fd_sc_hd__nand2_1
X_9432_ _7122_/X _6120_/Y _9475_/S vssd1 vssd1 vccd1 vccd1 _9432_/X sky130_fd_sc_hd__mux2_4
XFILLER_32_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6575_ _9676_/Q _6575_/B vssd1 vssd1 vccd1 vccd1 _6576_/B sky130_fd_sc_hd__or2_1
X_9363_ _7615_/X _7582_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9363_/X sky130_fd_sc_hd__mux2_1
X_5526_ _9380_/X _5505_/X _5611_/A vssd1 vssd1 vccd1 vccd1 _5605_/B sky130_fd_sc_hd__o21ai_1
X_9294_ _9293_/X input28/X _9294_/S vssd1 vssd1 vccd1 vccd1 _9294_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8314_ _4816_/X _8305_/Y _4814_/X _8111_/Y vssd1 vssd1 vccd1 vccd1 _8314_/X sky130_fd_sc_hd__o22a_1
XFILLER_132_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8245_ _6341_/A _8238_/B _8243_/Y vssd1 vssd1 vccd1 vccd1 _8245_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_117_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5457_ _9349_/X _9365_/X _5423_/Y _5491_/A vssd1 vssd1 vccd1 vccd1 _5457_/X sky130_fd_sc_hd__o22a_1
XFILLER_132_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8176_ _8176_/A _8998_/X vssd1 vssd1 vccd1 vccd1 _9522_/D sky130_fd_sc_hd__or2_1
X_5388_ _5388_/A vssd1 vssd1 vccd1 vccd1 _5389_/B sky130_fd_sc_hd__inv_2
XFILLER_59_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7127_ _7407_/A vssd1 vssd1 vccd1 vccd1 _7247_/A sky130_fd_sc_hd__buf_1
XFILLER_101_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7058_ _7058_/A vssd1 vssd1 vccd1 vccd1 _7079_/A sky130_fd_sc_hd__inv_2
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6009_ _6009_/A vssd1 vssd1 vccd1 vccd1 _6009_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6360_ _9751_/Q vssd1 vssd1 vccd1 vccd1 _6360_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5311_ _5222_/A _9732_/Q _5238_/B _5253_/Y vssd1 vssd1 vccd1 vccd1 _9732_/D sky130_fd_sc_hd__a22o_1
X_6291_ _9592_/Q _6171_/A _8042_/A _6142_/A vssd1 vssd1 vccd1 vccd1 _6296_/B sky130_fd_sc_hd__a22o_1
XFILLER_154_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8030_ _9460_/X _8030_/B vssd1 vssd1 vccd1 vccd1 _8030_/X sky130_fd_sc_hd__and2_1
XFILLER_5_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5242_ _5242_/A _5294_/A vssd1 vssd1 vccd1 vccd1 _5290_/A sky130_fd_sc_hd__or2_1
X_5173_ _9770_/Q _5167_/X input30/X _5168_/X _5165_/X vssd1 vssd1 vccd1 vccd1 _9770_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_110_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput1 io_QEI_ChA vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_1
XFILLER_68_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8932_ _8931_/A _8931_/B _8931_/X vssd1 vssd1 vccd1 vccd1 _8932_/X sky130_fd_sc_hd__a21bo_1
XFILLER_110_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8863_ _8863_/A _8862_/X vssd1 vssd1 vccd1 vccd1 _8863_/X sky130_fd_sc_hd__or2b_1
XFILLER_36_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7814_ _7814_/A _7814_/B vssd1 vssd1 vccd1 vccd1 _7819_/B sky130_fd_sc_hd__or2_1
XFILLER_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8794_ _8793_/A _8793_/B _8841_/A vssd1 vssd1 vccd1 vccd1 _8794_/X sky130_fd_sc_hd__a21bo_1
XFILLER_24_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7745_ _7743_/X _6353_/A _7797_/A _9753_/Q vssd1 vssd1 vccd1 vccd1 _7745_/X sky130_fd_sc_hd__o22a_1
X_4957_ _9113_/X _4951_/X _9850_/Q _4952_/X _4955_/X vssd1 vssd1 vccd1 vccd1 _9850_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7676_ _9919_/Q _7863_/A vssd1 vssd1 vccd1 vccd1 _7677_/B sky130_fd_sc_hd__or2_1
X_4888_ _9735_/Q _4865_/X _9883_/Q _4866_/X _4887_/X vssd1 vssd1 vccd1 vccd1 _9883_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9415_ _7124_/X _7492_/B _9475_/S vssd1 vssd1 vccd1 vccd1 _9415_/X sky130_fd_sc_hd__mux2_2
X_6627_ _6814_/A vssd1 vssd1 vccd1 vccd1 _6766_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_192_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6558_ _6558_/A _6558_/B vssd1 vssd1 vccd1 vccd1 _6575_/B sky130_fd_sc_hd__or2_1
X_9346_ _7058_/A _7610_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9346_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6489_ _6309_/Y _6475_/X _6478_/A _6480_/X vssd1 vssd1 vccd1 vccd1 _6489_/X sky130_fd_sc_hd__a211o_1
X_9277_ _9276_/X _7836_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9277_/X sky130_fd_sc_hd__mux2_1
X_5509_ _5507_/Y _5508_/Y _5507_/Y _5508_/Y vssd1 vssd1 vccd1 vccd1 _5509_/X sky130_fd_sc_hd__a2bb2o_4
X_8228_ _6429_/Y _8227_/Y _8225_/X vssd1 vssd1 vccd1 vccd1 _8228_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_120_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8159_ _7856_/A _8106_/X _8158_/X vssd1 vssd1 vccd1 vccd1 _8159_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5860_ _9627_/Q vssd1 vssd1 vccd1 vccd1 _5860_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4811_ _9286_/X _4809_/X _9913_/Q _4810_/X _4806_/X vssd1 vssd1 vccd1 vccd1 _9913_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5791_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5791_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4742_ _5136_/A vssd1 vssd1 vccd1 vccd1 _5128_/A sky130_fd_sc_hd__clkbuf_2
X_7530_ _7482_/A _7482_/B _7482_/X vssd1 vssd1 vccd1 vccd1 _7553_/A sky130_fd_sc_hd__a21bo_1
XFILLER_186_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7461_ _7459_/X _7460_/X _7459_/X _7460_/X vssd1 vssd1 vccd1 vccd1 _7461_/X sky130_fd_sc_hd__a2bb2o_2
X_9200_ _6544_/Y _9805_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9554_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6412_ _6347_/A _6390_/B _8203_/A vssd1 vssd1 vccd1 vccd1 _6416_/A sky130_fd_sc_hd__a21bo_1
XFILLER_147_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7392_ _7385_/A _7384_/B _7386_/A _7407_/B _7391_/Y vssd1 vssd1 vccd1 vccd1 _7393_/B
+ sky130_fd_sc_hd__o41a_1
X_6343_ _9777_/Q vssd1 vssd1 vccd1 vccd1 _6343_/Y sky130_fd_sc_hd__inv_2
X_9131_ _9868_/Q _9884_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9131_/X sky130_fd_sc_hd__mux2_1
X_6274_ _9589_/Q vssd1 vssd1 vccd1 vccd1 _8036_/A sky130_fd_sc_hd__inv_2
XFILLER_170_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9062_ _8032_/Y _8031_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9062_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8013_ _8013_/A _8021_/B vssd1 vssd1 vccd1 vccd1 _8013_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5225_ _9745_/Q vssd1 vssd1 vccd1 vccd1 _5250_/A sky130_fd_sc_hd__inv_2
XFILLER_130_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5156_ _5179_/A vssd1 vssd1 vccd1 vccd1 _5205_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5087_ _5084_/X _6318_/A _5086_/Y _5073_/X vssd1 vssd1 vccd1 vccd1 _5088_/B sky130_fd_sc_hd__o22a_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8915_ _8907_/X _8914_/X _8907_/X _8914_/X vssd1 vssd1 vccd1 vccd1 _8915_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_25_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9895_ _9895_/CLK _9895_/D vssd1 vssd1 vccd1 vccd1 _9895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8846_ _8845_/A _8845_/B _8944_/A vssd1 vssd1 vccd1 vccd1 _8846_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_112_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8777_ _5852_/X _8656_/X _8776_/X vssd1 vssd1 vccd1 vccd1 _8777_/Y sky130_fd_sc_hd__a21oi_1
X_5989_ _5989_/A _5989_/B vssd1 vssd1 vccd1 vccd1 _5989_/X sky130_fd_sc_hd__or2_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7728_ _7873_/A vssd1 vssd1 vccd1 vccd1 _7728_/X sky130_fd_sc_hd__buf_2
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7659_ _9902_/Q _7659_/B vssd1 vssd1 vccd1 vccd1 _7795_/A sky130_fd_sc_hd__or2_1
XFILLER_20_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9329_ _9328_/X _7907_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9329_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5010_ _9829_/Q _5003_/X input24/X _5004_/X _5008_/X vssd1 vssd1 vccd1 vccd1 _9829_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_112_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_clock/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8700_ _8699_/A _8699_/B _8747_/A vssd1 vssd1 vccd1 vccd1 _8700_/X sky130_fd_sc_hd__a21o_1
X_6961_ _6909_/X _6912_/X _6913_/X _6960_/X vssd1 vssd1 vccd1 vccd1 _6964_/A sky130_fd_sc_hd__o22a_1
XFILLER_81_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9680_ _9699_/CLK _9680_/D vssd1 vssd1 vccd1 vccd1 _9680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5912_ _5915_/A _9131_/X vssd1 vssd1 vccd1 vccd1 _9599_/D sky130_fd_sc_hd__and2_1
X_6892_ _6892_/A vssd1 vssd1 vccd1 vccd1 _6892_/Y sky130_fd_sc_hd__inv_2
X_8631_ _8629_/Y _8630_/X _8629_/Y _8630_/X vssd1 vssd1 vccd1 vccd1 _8631_/X sky130_fd_sc_hd__o2bb2a_1
X_5843_ _9634_/Q vssd1 vssd1 vccd1 vccd1 _5843_/X sky130_fd_sc_hd__buf_2
XFILLER_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8562_ _8534_/A _9382_/X _8472_/A _8773_/B vssd1 vssd1 vccd1 vccd1 _8564_/A sky130_fd_sc_hd__o22a_1
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5774_ _8967_/B vssd1 vssd1 vccd1 vccd1 _5774_/X sky130_fd_sc_hd__clkbuf_2
X_7513_ _7202_/X _7511_/X _7145_/A _7512_/X vssd1 vssd1 vccd1 vccd1 _7514_/B sky130_fd_sc_hd__o22a_1
XFILLER_21_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8493_ _9382_/X vssd1 vssd1 vccd1 vccd1 _8652_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7444_ _7441_/X _7443_/X _7441_/X _7443_/X vssd1 vssd1 vccd1 vccd1 _7444_/X sky130_fd_sc_hd__a2bb2o_1
X_7375_ _7298_/A _7304_/A _7298_/Y vssd1 vssd1 vccd1 vccd1 _7376_/B sky130_fd_sc_hd__a21o_1
X_6326_ _8186_/A vssd1 vssd1 vccd1 vccd1 _8056_/A sky130_fd_sc_hd__clkbuf_2
X_9114_ _9598_/Q _5035_/A _9667_/Q vssd1 vssd1 vccd1 vccd1 _9114_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6257_ _6265_/A _6265_/B _6248_/Y _6256_/X vssd1 vssd1 vccd1 vccd1 _6257_/X sky130_fd_sc_hd__o31a_1
X_9045_ _8001_/Y _9608_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9045_/X sky130_fd_sc_hd__mux2_1
X_5208_ _5026_/X _5203_/X _9755_/Q _5205_/X _5206_/X vssd1 vssd1 vccd1 vccd1 _9755_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6188_ _7976_/A _6137_/A _7983_/A _6137_/A vssd1 vssd1 vccd1 vccd1 _6189_/B sky130_fd_sc_hd__o22a_1
X_5139_ _5136_/X _9785_/Q _5138_/X _9212_/X _5132_/X vssd1 vssd1 vccd1 vccd1 _9785_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_123_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9878_ _9879_/CLK _9878_/D vssd1 vssd1 vccd1 vccd1 _9878_/Q sky130_fd_sc_hd__dfxtp_1
X_8829_ _8829_/A _8959_/B _8734_/X vssd1 vssd1 vccd1 vccd1 _8829_/X sky130_fd_sc_hd__or3b_1
XFILLER_80_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_6_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _9836_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5490_ _9476_/X _5489_/X _9476_/X _5489_/X vssd1 vssd1 vccd1 vccd1 _5588_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7160_ _7160_/A _9431_/X vssd1 vssd1 vccd1 vccd1 _7548_/A sky130_fd_sc_hd__or2_1
XFILLER_98_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6111_ _9863_/Q _9650_/Q _8008_/A _6110_/Y vssd1 vssd1 vccd1 vccd1 _6111_/X sky130_fd_sc_hd__o22a_1
XFILLER_98_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7091_ _7088_/A _7088_/B _7089_/B vssd1 vssd1 vccd1 vccd1 _7091_/X sky130_fd_sc_hd__a21bo_1
X_6042_ _9856_/Q vssd1 vssd1 vccd1 vccd1 _7974_/A sky130_fd_sc_hd__inv_2
XFILLER_39_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9801_ _9923_/CLK _9801_/D vssd1 vssd1 vccd1 vccd1 _9801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7993_ _7993_/A _7993_/B vssd1 vssd1 vccd1 vccd1 _7993_/Y sky130_fd_sc_hd__nor2_1
X_9732_ _9893_/CLK _9732_/D vssd1 vssd1 vccd1 vccd1 _9732_/Q sky130_fd_sc_hd__dfxtp_1
X_6944_ _6902_/A _6902_/B _6903_/B vssd1 vssd1 vccd1 vccd1 _6944_/X sky130_fd_sc_hd__a21bo_1
X_9663_ _9673_/CLK _9663_/D vssd1 vssd1 vccd1 vccd1 _9663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8614_ _8614_/A vssd1 vssd1 vccd1 vccd1 _8614_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6875_ _6868_/A _6867_/B _6867_/C _6877_/A _6874_/Y vssd1 vssd1 vccd1 vccd1 _6876_/B
+ sky130_fd_sc_hd__o41a_1
XFILLER_22_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9594_ _9924_/CLK _9594_/D vssd1 vssd1 vccd1 vccd1 _9594_/Q sky130_fd_sc_hd__dfxtp_1
X_5826_ _9647_/Q _5824_/X input19/X _5825_/X _5822_/X vssd1 vssd1 vccd1 vccd1 _9647_/D
+ sky130_fd_sc_hd__o221a_1
X_8545_ _8630_/A _9379_/X _8545_/C vssd1 vssd1 vccd1 vccd1 _8547_/A sky130_fd_sc_hd__or3_4
X_5757_ _6598_/A _5713_/Y _5714_/X _5756_/X vssd1 vssd1 vccd1 vccd1 _5757_/Y sky130_fd_sc_hd__o22ai_4
X_8476_ _8455_/Y _8475_/X _8455_/Y _8475_/X vssd1 vssd1 vccd1 vccd1 _8476_/X sky130_fd_sc_hd__o2bb2a_2
XFILLER_182_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5688_ _8389_/B _5681_/X _9102_/X _5684_/X _5682_/X vssd1 vssd1 vccd1 vccd1 _9675_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_108_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7427_ _7427_/A _7427_/B vssd1 vssd1 vccd1 vccd1 _7428_/B sky130_fd_sc_hd__nor2_1
XFILLER_162_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7358_ _7356_/X _7357_/X _7356_/X _7357_/X vssd1 vssd1 vccd1 vccd1 _7358_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_150_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6309_ _9784_/Q vssd1 vssd1 vccd1 vccd1 _6309_/Y sky130_fd_sc_hd__inv_2
X_7289_ _7276_/X _7277_/X _7276_/X _7277_/X vssd1 vssd1 vccd1 vccd1 _7289_/X sky130_fd_sc_hd__a2bb2o_2
X_9028_ _9027_/X _9755_/Q _9481_/S vssd1 vssd1 vccd1 vccd1 _9028_/X sky130_fd_sc_hd__mux2_2
XFILLER_49_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4990_ _9841_/Q _4985_/X input37/X _4987_/X _4974_/X vssd1 vssd1 vccd1 vccd1 _9841_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6660_ _6660_/A _6660_/B vssd1 vssd1 vccd1 vccd1 _6672_/A sky130_fd_sc_hd__or2_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5611_ _5611_/A vssd1 vssd1 vccd1 vccd1 _5611_/Y sky130_fd_sc_hd__inv_2
X_6591_ _8381_/B vssd1 vssd1 vccd1 vccd1 _6591_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5542_ _9384_/X _5477_/X _5565_/A vssd1 vssd1 vccd1 vccd1 _5561_/B sky130_fd_sc_hd__o21ai_1
X_8330_ _7665_/A _8308_/Y _4820_/X _8306_/Y _8311_/X vssd1 vssd1 vccd1 vccd1 _8330_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_191_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8261_ _8189_/X _8260_/X _8189_/X _8260_/X vssd1 vssd1 vccd1 vccd1 _8261_/X sky130_fd_sc_hd__o2bb2a_1
X_5473_ _5471_/Y _5472_/Y _5471_/Y _5472_/Y vssd1 vssd1 vccd1 vccd1 _5473_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_172_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8192_ _8235_/B vssd1 vssd1 vccd1 vccd1 _8231_/B sky130_fd_sc_hd__buf_2
X_7212_ _9626_/Q vssd1 vssd1 vccd1 vccd1 _7384_/C sky130_fd_sc_hd__inv_2
X_7143_ _9430_/X vssd1 vssd1 vccd1 vccd1 _7522_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_113_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7074_ _7074_/A _7074_/B vssd1 vssd1 vccd1 vccd1 _7075_/B sky130_fd_sc_hd__or2_1
XFILLER_58_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6025_ _9854_/Q _6023_/Y _7962_/A _9641_/Q vssd1 vssd1 vccd1 vccd1 _6026_/A sky130_fd_sc_hd__o22a_2
XFILLER_104_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9715_ _9715_/CLK _9715_/D vssd1 vssd1 vccd1 vccd1 _9715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7976_ _7976_/A _7993_/B vssd1 vssd1 vccd1 vccd1 _7976_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6927_ _6924_/X _6926_/X _6924_/X _6926_/X vssd1 vssd1 vccd1 vccd1 _6927_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9646_ _9650_/CLK _9646_/D vssd1 vssd1 vccd1 vccd1 _9646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6858_ _6781_/A _6787_/A _6781_/Y vssd1 vssd1 vccd1 vccd1 _6859_/B sky130_fd_sc_hd__a21o_1
XFILLER_196_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5809_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5809_/X sky130_fd_sc_hd__buf_2
XFILLER_13_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9577_ _9578_/CLK _9577_/D vssd1 vssd1 vccd1 vccd1 _9577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8528_ _8499_/Y _8504_/X _8505_/X _8506_/Y vssd1 vssd1 vccd1 vccd1 _8528_/X sky130_fd_sc_hd__o22a_1
X_6789_ _6767_/X _6788_/X _6767_/X _6788_/X vssd1 vssd1 vccd1 vccd1 _6789_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8459_ _8457_/A _8457_/B _8478_/A vssd1 vssd1 vccd1 vccd1 _8460_/B sky130_fd_sc_hd__a21o_1
XFILLER_163_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_24_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _9715_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_39_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _9910_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7830_ _4816_/X _7667_/B _7829_/Y vssd1 vssd1 vccd1 vccd1 _7830_/X sky130_fd_sc_hd__a21o_1
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4973_ _9846_/Q vssd1 vssd1 vccd1 vccd1 _4973_/X sky130_fd_sc_hd__buf_2
X_7761_ _7827_/A vssd1 vssd1 vccd1 vccd1 _7761_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7692_ _7856_/A vssd1 vssd1 vccd1 vccd1 _7692_/X sky130_fd_sc_hd__clkbuf_2
X_9500_ _9499_/X _8919_/A _9505_/S vssd1 vssd1 vccd1 vccd1 _9500_/X sky130_fd_sc_hd__mux2_1
X_6712_ _6868_/A _6842_/A vssd1 vssd1 vccd1 vccd1 _6713_/C sky130_fd_sc_hd__or2_2
XFILLER_32_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6643_ _6756_/A _6691_/B _7030_/A vssd1 vssd1 vccd1 vccd1 _6644_/B sky130_fd_sc_hd__and3_1
X_9431_ _7119_/X _5785_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9431_/X sky130_fd_sc_hd__mux2_2
XFILLER_32_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6574_ _6571_/Y _6573_/X _6553_/B vssd1 vssd1 vccd1 vccd1 _6574_/Y sky130_fd_sc_hd__o21ai_1
X_9362_ _7065_/A _7624_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9362_/X sky130_fd_sc_hd__mux2_1
X_5525_ _5612_/A _5612_/B vssd1 vssd1 vccd1 vccd1 _5611_/A sky130_fd_sc_hd__nand2_1
X_9293_ _9292_/X _7862_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9293_/X sky130_fd_sc_hd__mux2_1
X_8313_ _7665_/A _8308_/Y _4820_/X _8306_/Y _8312_/Y vssd1 vssd1 vccd1 vccd1 _8313_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_160_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8244_ _6339_/Y _8243_/Y _8240_/B vssd1 vssd1 vccd1 vccd1 _8244_/Y sky130_fd_sc_hd__o21ai_1
X_5456_ _9357_/X _9355_/X _5426_/Y _5495_/A vssd1 vssd1 vccd1 vccd1 _5491_/A sky130_fd_sc_hd__o22a_1
XFILLER_160_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8175_ _8175_/A _8174_/X vssd1 vssd1 vccd1 vccd1 _9562_/D sky130_fd_sc_hd__nor2b_1
X_5387_ _5387_/A vssd1 vssd1 vccd1 vccd1 _9721_/D sky130_fd_sc_hd__inv_2
XFILLER_101_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7126_ _7384_/A vssd1 vssd1 vccd1 vccd1 _7407_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7057_ _7057_/A vssd1 vssd1 vccd1 vccd1 _7080_/A sky130_fd_sc_hd__inv_2
X_6008_ _6008_/A _6008_/B vssd1 vssd1 vccd1 vccd1 _6009_/A sky130_fd_sc_hd__or2_1
XFILLER_86_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7959_ _8543_/A vssd1 vssd1 vccd1 vccd1 _8773_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_131_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9629_ _9634_/CLK _9629_/D vssd1 vssd1 vccd1 vccd1 _9629_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6290_ _9592_/Q vssd1 vssd1 vccd1 vccd1 _8042_/A sky130_fd_sc_hd__inv_2
XFILLER_154_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5310_ _5310_/A vssd1 vssd1 vccd1 vccd1 _9733_/D sky130_fd_sc_hd__inv_2
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5241_ _5241_/A _5298_/A vssd1 vssd1 vccd1 vccd1 _5294_/A sky130_fd_sc_hd__or2_1
X_5172_ _9771_/Q _5167_/X input31/X _5168_/X _5165_/X vssd1 vssd1 vccd1 vccd1 _9771_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_122_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput2 io_QEI_ChB vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
X_8931_ _8931_/A _8931_/B vssd1 vssd1 vccd1 vccd1 _8931_/X sky130_fd_sc_hd__or2_1
XFILLER_110_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8862_ _8944_/C _9422_/X _8935_/A _9429_/X vssd1 vssd1 vccd1 vccd1 _8862_/X sky130_fd_sc_hd__or4_4
X_8793_ _8793_/A _8793_/B vssd1 vssd1 vccd1 vccd1 _8841_/A sky130_fd_sc_hd__or2_1
X_7813_ _9906_/Q _7663_/B _7812_/Y vssd1 vssd1 vccd1 vccd1 _7813_/X sky130_fd_sc_hd__a21o_1
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7744_ _9902_/Q vssd1 vssd1 vccd1 vccd1 _7797_/A sky130_fd_sc_hd__inv_2
XFILLER_24_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4956_ _9114_/X _4951_/X _9851_/Q _4952_/X _4955_/X vssd1 vssd1 vccd1 vccd1 _9851_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7675_ _9918_/Q _7675_/B vssd1 vssd1 vccd1 vccd1 _7863_/A sky130_fd_sc_hd__or2_1
X_4887_ _5206_/A vssd1 vssd1 vccd1 vccd1 _4887_/X sky130_fd_sc_hd__buf_2
XFILLER_51_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9414_ _7123_/X _6119_/Y _9475_/S vssd1 vssd1 vccd1 vccd1 _9414_/X sky130_fd_sc_hd__mux2_2
X_6626_ _6796_/D vssd1 vssd1 vccd1 vccd1 _6814_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_192_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6557_ _6561_/A _6557_/B vssd1 vssd1 vccd1 vccd1 _6558_/B sky130_fd_sc_hd__or2_1
X_9345_ _7069_/A _7630_/Y _9683_/Q vssd1 vssd1 vccd1 vccd1 _9345_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5508_ _5434_/A _5434_/B _5434_/Y vssd1 vssd1 vccd1 vccd1 _5508_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_173_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6488_ _6485_/X _6486_/X _6487_/X vssd1 vssd1 vccd1 vccd1 _6488_/X sky130_fd_sc_hd__a21o_1
X_9276_ _9762_/Q _9275_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9276_/X sky130_fd_sc_hd__mux2_1
X_8227_ _8227_/A _8227_/B vssd1 vssd1 vccd1 vccd1 _8227_/Y sky130_fd_sc_hd__nor2_2
XFILLER_79_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5439_ _9668_/Q vssd1 vssd1 vccd1 vccd1 _5442_/A sky130_fd_sc_hd__inv_2
XFILLER_126_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8158_ _7738_/A _8107_/X _8157_/X vssd1 vssd1 vccd1 vccd1 _8158_/X sky130_fd_sc_hd__a21o_1
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7109_ _7109_/A _7109_/B vssd1 vssd1 vccd1 vccd1 _7110_/B sky130_fd_sc_hd__or2_1
X_8089_ _9559_/Q _8089_/B vssd1 vssd1 vccd1 vccd1 _8089_/X sky130_fd_sc_hd__or2_1
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4810_ _4836_/A vssd1 vssd1 vccd1 vccd1 _4810_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5790_ _5790_/A vssd1 vssd1 vccd1 vccd1 _5840_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4741_ _9929_/Q vssd1 vssd1 vccd1 vccd1 _5136_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_202_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7460_ _7358_/X _7369_/X _7358_/X _7369_/X vssd1 vssd1 vccd1 vccd1 _7460_/X sky130_fd_sc_hd__a2bb2o_2
X_6411_ _6544_/B vssd1 vssd1 vccd1 vccd1 _6411_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9130_ _9867_/Q _9883_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9130_/X sky130_fd_sc_hd__mux2_1
X_7391_ _7394_/C _7391_/B vssd1 vssd1 vccd1 vccd1 _7391_/Y sky130_fd_sc_hd__nand2_1
X_6342_ _9778_/Q vssd1 vssd1 vccd1 vccd1 _6342_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6273_ _6271_/X _6272_/Y _6271_/X _6272_/Y vssd1 vssd1 vccd1 vccd1 _6273_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_170_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9061_ _8030_/X _8029_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9061_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8012_ _8046_/B vssd1 vssd1 vccd1 vccd1 _8021_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_102_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5224_ _5224_/A vssd1 vssd1 vccd1 vccd1 _5224_/X sky130_fd_sc_hd__clkbuf_2
X_5155_ _5178_/A vssd1 vssd1 vccd1 vccd1 _5155_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5086_ _9835_/Q vssd1 vssd1 vccd1 vccd1 _5086_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8914_ _8913_/A _8913_/B _8913_/Y vssd1 vssd1 vccd1 vccd1 _8914_/X sky130_fd_sc_hd__a21o_1
X_9894_ _9895_/CLK _9894_/D vssd1 vssd1 vccd1 vccd1 _9894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8845_ _8845_/A _8845_/B vssd1 vssd1 vccd1 vccd1 _8944_/A sky130_fd_sc_hd__nand2_1
XFILLER_112_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8776_ _8776_/A _8800_/B vssd1 vssd1 vccd1 vccd1 _8776_/X sky130_fd_sc_hd__or2_1
X_5988_ _9849_/Q _5979_/Y _5704_/B _5981_/Y vssd1 vssd1 vccd1 vccd1 _5989_/B sky130_fd_sc_hd__o22a_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7727_ _9920_/Q vssd1 vssd1 vccd1 vccd1 _7873_/A sky130_fd_sc_hd__inv_2
XFILLER_12_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4939_ _4991_/A vssd1 vssd1 vccd1 vccd1 _4939_/X sky130_fd_sc_hd__buf_1
X_7658_ _7793_/A _7658_/B vssd1 vssd1 vccd1 vccd1 _7659_/B sky130_fd_sc_hd__nand2_1
XFILLER_138_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6609_ _6660_/B vssd1 vssd1 vccd1 vccd1 _7005_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_137_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7589_ _7589_/A vssd1 vssd1 vccd1 vccd1 _7593_/A sky130_fd_sc_hd__inv_2
X_9328_ _9778_/Q _9327_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9328_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9259_ _7813_/X _9757_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9259_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6960_ _6914_/X _6919_/X _6920_/X _6959_/X vssd1 vssd1 vccd1 vccd1 _6960_/X sky130_fd_sc_hd__o22a_1
X_5911_ _5915_/A _9132_/X vssd1 vssd1 vccd1 vccd1 _9600_/D sky130_fd_sc_hd__and2_1
XFILLER_179_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6891_ _9618_/Q _6891_/B _6902_/A vssd1 vssd1 vccd1 vccd1 _6892_/A sky130_fd_sc_hd__and3_1
X_8630_ _8630_/A _8766_/B _8630_/C vssd1 vssd1 vccd1 vccd1 _8630_/X sky130_fd_sc_hd__or3_1
X_5842_ _9635_/Q _5832_/A _5041_/X _5833_/A _5840_/X vssd1 vssd1 vccd1 vccd1 _9635_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8561_ _8533_/X _8539_/X _8540_/X _8541_/X vssd1 vssd1 vccd1 vccd1 _8561_/X sky130_fd_sc_hd__o22a_1
X_5773_ _9663_/Q _5697_/X _5769_/X _7120_/A _5772_/X vssd1 vssd1 vccd1 vccd1 _9663_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_147_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7512_ _7202_/X _7511_/X _7202_/X _7511_/X vssd1 vssd1 vccd1 vccd1 _7512_/X sky130_fd_sc_hd__a2bb2o_1
X_8492_ _8491_/A _8491_/B _8526_/A vssd1 vssd1 vccd1 vccd1 _8492_/X sky130_fd_sc_hd__a21bo_1
X_7443_ _7443_/A _7443_/B vssd1 vssd1 vccd1 vccd1 _7443_/X sky130_fd_sc_hd__or2_1
XFILLER_174_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7374_ _7374_/A _7374_/B vssd1 vssd1 vccd1 vccd1 _7376_/A sky130_fd_sc_hd__or2_1
X_6325_ _9844_/Q vssd1 vssd1 vccd1 vccd1 _8186_/A sky130_fd_sc_hd__inv_2
XFILLER_115_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9113_ _9597_/Q _4860_/A _9667_/Q vssd1 vssd1 vccd1 vccd1 _9113_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9044_ _7998_/Y _9043_/X _9053_/S vssd1 vssd1 vccd1 vccd1 _9044_/X sky130_fd_sc_hd__mux2_1
X_6256_ _8021_/A _6245_/X _8024_/A _6245_/X vssd1 vssd1 vccd1 vccd1 _6256_/X sky130_fd_sc_hd__o22a_1
X_5207_ input46/X _5203_/X _6341_/A _5205_/X _5206_/X vssd1 vssd1 vccd1 vccd1 _9756_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6187_ _6187_/A _6187_/B vssd1 vssd1 vccd1 vccd1 _6200_/C sky130_fd_sc_hd__or2_1
X_5138_ _5138_/A vssd1 vssd1 vccd1 vccd1 _5138_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5069_ _5069_/A _5069_/B vssd1 vssd1 vccd1 vccd1 _9807_/D sky130_fd_sc_hd__nor2_1
X_9877_ _9879_/CLK _9877_/D vssd1 vssd1 vccd1 vccd1 _9877_/Q sky130_fd_sc_hd__dfxtp_1
X_8828_ _9396_/X vssd1 vssd1 vccd1 vccd1 _8959_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_25_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8759_ _8757_/X _8826_/A _8757_/X _8826_/A vssd1 vssd1 vccd1 vccd1 _8760_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_181_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6110_ _9650_/Q vssd1 vssd1 vccd1 vccd1 _6110_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7090_ _7089_/A _7089_/B _7107_/B vssd1 vssd1 vccd1 vccd1 _7090_/X sky130_fd_sc_hd__a21bo_1
X_6041_ _9643_/Q vssd1 vssd1 vccd1 vccd1 _6041_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9800_ _9833_/CLK _9800_/D vssd1 vssd1 vccd1 vccd1 _9800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7992_ _8990_/X _8009_/B vssd1 vssd1 vccd1 vccd1 _7992_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9731_ _9879_/CLK _9731_/D vssd1 vssd1 vccd1 vccd1 _9731_/Q sky130_fd_sc_hd__dfxtp_1
X_6943_ _6841_/X _6852_/X _6841_/X _6852_/X vssd1 vssd1 vccd1 vccd1 _6943_/X sky130_fd_sc_hd__a2bb2o_1
X_9662_ _9673_/CLK _9662_/D vssd1 vssd1 vccd1 vccd1 _9662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6874_ _6877_/C _6874_/B vssd1 vssd1 vccd1 vccd1 _6874_/Y sky130_fd_sc_hd__nand2_1
X_8613_ _8613_/A _8568_/X vssd1 vssd1 vccd1 vccd1 _8614_/A sky130_fd_sc_hd__or2b_1
X_5825_ _5833_/A vssd1 vssd1 vccd1 vccd1 _5825_/X sky130_fd_sc_hd__clkbuf_2
X_9593_ _9924_/CLK _9593_/D vssd1 vssd1 vccd1 vccd1 _9593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8544_ _8606_/A _8625_/B vssd1 vssd1 vccd1 vccd1 _8546_/A sky130_fd_sc_hd__or2_2
X_5756_ _8381_/B _9664_/Q _5715_/Y _5755_/X vssd1 vssd1 vccd1 vccd1 _5756_/X sky130_fd_sc_hd__o2bb2a_1
X_8475_ _8475_/A _8584_/B _8475_/C vssd1 vssd1 vccd1 vccd1 _8475_/X sky130_fd_sc_hd__or3_1
XFILLER_163_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5687_ _9676_/Q _5681_/X _9103_/X _5684_/X _5682_/X vssd1 vssd1 vccd1 vccd1 _9676_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_175_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7426_ _7378_/X _7423_/X _7424_/X _7425_/X vssd1 vssd1 vccd1 vccd1 _7426_/X sky130_fd_sc_hd__o22a_1
XFILLER_162_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7357_ _7302_/A _7302_/B _7303_/B vssd1 vssd1 vccd1 vccd1 _7357_/X sky130_fd_sc_hd__a21bo_1
X_6308_ _4973_/X _6304_/Y _4976_/X _6487_/A _6307_/X vssd1 vssd1 vccd1 vccd1 _6308_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_143_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7288_ _7288_/A _7288_/B vssd1 vssd1 vccd1 vccd1 _7299_/A sky130_fd_sc_hd__or2_2
X_9027_ _9787_/Q _9904_/Q _9480_/S vssd1 vssd1 vccd1 vccd1 _9027_/X sky130_fd_sc_hd__mux2_1
X_6239_ _6244_/B _6238_/Y _6244_/B _6238_/Y vssd1 vssd1 vccd1 vccd1 _6239_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9929_ _9929_/CLK _9929_/D vssd1 vssd1 vccd1 vccd1 _9929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5610_ _8177_/A vssd1 vssd1 vccd1 vccd1 _8176_/A sky130_fd_sc_hd__buf_2
X_6590_ _6660_/A vssd1 vssd1 vccd1 vccd1 _6975_/A sky130_fd_sc_hd__buf_2
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5541_ _5566_/A _5566_/B vssd1 vssd1 vccd1 vccd1 _5565_/A sky130_fd_sc_hd__or2_1
XFILLER_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8260_ _8051_/A _8183_/B _8183_/Y vssd1 vssd1 vccd1 vccd1 _8260_/X sky130_fd_sc_hd__a21o_1
XFILLER_129_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5472_ _5409_/A _5409_/B _5409_/Y vssd1 vssd1 vccd1 vccd1 _5472_/Y sky130_fd_sc_hd__a21oi_1
X_7211_ _9469_/X vssd1 vssd1 vccd1 vccd1 _7283_/B sky130_fd_sc_hd__clkbuf_2
X_8191_ _8191_/A _8191_/B vssd1 vssd1 vccd1 vccd1 _8235_/B sky130_fd_sc_hd__nand2_1
XFILLER_144_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7142_ _7394_/A vssd1 vssd1 vccd1 vccd1 _7234_/A sky130_fd_sc_hd__buf_2
X_7073_ _7073_/A _7073_/B vssd1 vssd1 vccd1 vccd1 _7074_/B sky130_fd_sc_hd__or2_1
XFILLER_58_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6024_ _9854_/Q vssd1 vssd1 vccd1 vccd1 _7962_/A sky130_fd_sc_hd__inv_2
XFILLER_100_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_5_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _9923_/CLK sky130_fd_sc_hd__clkbuf_16
X_7975_ _9371_/X _7987_/B vssd1 vssd1 vccd1 vccd1 _7975_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9714_ _9828_/CLK _9714_/D vssd1 vssd1 vccd1 vccd1 _9714_/Q sky130_fd_sc_hd__dfxtp_1
X_6926_ _6926_/A _6926_/B vssd1 vssd1 vccd1 vccd1 _6926_/X sky130_fd_sc_hd__or2_1
XFILLER_54_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9645_ _9828_/CLK _9645_/D vssd1 vssd1 vccd1 vccd1 _9645_/Q sky130_fd_sc_hd__dfxtp_2
X_6857_ _6857_/A _6857_/B vssd1 vssd1 vccd1 vccd1 _6859_/A sky130_fd_sc_hd__or2_1
XFILLER_210_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5808_ _5808_/A vssd1 vssd1 vccd1 vccd1 _7084_/A sky130_fd_sc_hd__inv_2
X_9576_ _9910_/CLK _9576_/D vssd1 vssd1 vccd1 vccd1 _9576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6788_ _6782_/A _6777_/X _6781_/Y _6779_/A _6787_/Y vssd1 vssd1 vccd1 vccd1 _6788_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_195_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8527_ _8526_/A _8526_/B _8559_/A vssd1 vssd1 vccd1 vccd1 _8527_/X sky130_fd_sc_hd__a21o_1
X_5739_ _9672_/Q _9655_/Q _6564_/A _5738_/Y vssd1 vssd1 vccd1 vccd1 _5739_/X sky130_fd_sc_hd__a22o_1
XFILLER_10_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8458_ _8458_/A vssd1 vssd1 vccd1 vccd1 _8478_/A sky130_fd_sc_hd__inv_2
XFILLER_175_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8389_ _8389_/A _8389_/B vssd1 vssd1 vccd1 vccd1 _8389_/Y sky130_fd_sc_hd__nor2_1
X_7409_ _7409_/A vssd1 vssd1 vccd1 vccd1 _7409_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4972_ _4969_/A _4969_/B _4969_/Y vssd1 vssd1 vccd1 vccd1 _4972_/Y sky130_fd_sc_hd__a21oi_1
X_7760_ _9909_/Q vssd1 vssd1 vccd1 vccd1 _7827_/A sky130_fd_sc_hd__inv_2
XFILLER_63_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7691_ _9916_/Q vssd1 vssd1 vccd1 vccd1 _7856_/A sky130_fd_sc_hd__inv_2
X_6711_ _6756_/B vssd1 vssd1 vccd1 vccd1 _6774_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_177_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6642_ _6642_/A _9464_/X vssd1 vssd1 vccd1 vccd1 _7030_/A sky130_fd_sc_hd__or2_2
X_9430_ _7118_/X _5782_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9430_/X sky130_fd_sc_hd__mux2_4
XFILLER_32_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9361_ _7060_/A _7614_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9361_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6573_ _6890_/A vssd1 vssd1 vccd1 vccd1 _6573_/X sky130_fd_sc_hd__buf_2
X_8312_ _8328_/B _8310_/X _8311_/X vssd1 vssd1 vccd1 vccd1 _8312_/Y sky130_fd_sc_hd__o21ai_1
X_5524_ _9446_/X _5509_/X _5616_/A vssd1 vssd1 vccd1 vccd1 _5612_/B sky130_fd_sc_hd__o21ai_1
X_9292_ _9768_/Q _9291_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9292_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8243_ _8243_/A vssd1 vssd1 vccd1 vccd1 _8243_/Y sky130_fd_sc_hd__inv_2
X_5455_ _9364_/X _9362_/X _5427_/X _5454_/X vssd1 vssd1 vccd1 vccd1 _5495_/A sky130_fd_sc_hd__o22a_1
X_8174_ _8174_/A _8174_/B vssd1 vssd1 vccd1 vccd1 _8174_/X sky130_fd_sc_hd__or2_1
XFILLER_117_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5386_ _5381_/B _5379_/X _5385_/Y _5328_/A _5364_/A vssd1 vssd1 vccd1 vccd1 _5387_/A
+ sky130_fd_sc_hd__o32a_1
X_7125_ _9625_/Q vssd1 vssd1 vccd1 vccd1 _7384_/A sky130_fd_sc_hd__inv_2
XFILLER_113_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7056_ _7056_/A vssd1 vssd1 vccd1 vccd1 _7081_/A sky130_fd_sc_hd__inv_2
X_6007_ _5989_/X _5998_/A _6006_/X vssd1 vssd1 vccd1 vccd1 _6008_/B sky130_fd_sc_hd__o21ba_1
XFILLER_86_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7958_ _9633_/Q vssd1 vssd1 vccd1 vccd1 _8543_/A sky130_fd_sc_hd__inv_2
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7889_ _7889_/A vssd1 vssd1 vccd1 vccd1 _7889_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6909_ _6861_/X _6906_/X _6907_/X _6908_/X vssd1 vssd1 vccd1 vccd1 _6909_/X sky130_fd_sc_hd__o22a_1
XFILLER_42_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9628_ _9634_/CLK _9628_/D vssd1 vssd1 vccd1 vccd1 _9628_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9559_ _9928_/CLK _9559_/D vssd1 vssd1 vccd1 vccd1 _9559_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240_ _5240_/A _5305_/A _5240_/C vssd1 vssd1 vccd1 vccd1 _5298_/A sky130_fd_sc_hd__or3_1
XFILLER_130_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5171_ _6347_/A _5167_/X input32/X _5168_/X _5165_/X vssd1 vssd1 vccd1 vccd1 _9772_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_122_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8930_ _8930_/A vssd1 vssd1 vccd1 vccd1 _8931_/B sky130_fd_sc_hd__inv_2
Xinput3 io_wb_adr_i[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_4
X_8861_ _8755_/A _9422_/X _8829_/A _8942_/B vssd1 vssd1 vccd1 vccd1 _8863_/A sky130_fd_sc_hd__o22a_1
X_8792_ _8792_/A vssd1 vssd1 vccd1 vccd1 _8793_/B sky130_fd_sc_hd__inv_2
X_7812_ _7812_/A vssd1 vssd1 vccd1 vccd1 _7812_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4955_ _4991_/A vssd1 vssd1 vccd1 vccd1 _4955_/X sky130_fd_sc_hd__buf_2
X_7743_ _7743_/A vssd1 vssd1 vccd1 vccd1 _7743_/X sky130_fd_sc_hd__buf_2
XFILLER_51_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7674_ _9917_/Q _7854_/A vssd1 vssd1 vccd1 vccd1 _7675_/B sky130_fd_sc_hd__or2_1
X_4886_ _9736_/Q _4879_/X _9884_/Q _4880_/X _4881_/X vssd1 vssd1 vccd1 vccd1 _9884_/D
+ sky130_fd_sc_hd__a221o_1
X_9413_ _9412_/X _7005_/A _9507_/S vssd1 vssd1 vccd1 vccd1 _9413_/X sky130_fd_sc_hd__mux2_1
X_6625_ _9614_/Q vssd1 vssd1 vccd1 vccd1 _6796_/D sky130_fd_sc_hd__inv_2
XFILLER_192_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6556_ _6556_/A _6556_/B vssd1 vssd1 vccd1 vccd1 _6557_/B sky130_fd_sc_hd__or2_1
X_9344_ _7609_/X _7564_/Y _9475_/S vssd1 vssd1 vccd1 vccd1 _9344_/X sky130_fd_sc_hd__mux2_4
XFILLER_192_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9275_ _7834_/Y _9762_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9275_/X sky130_fd_sc_hd__mux2_1
X_5507_ _5507_/A vssd1 vssd1 vccd1 vccd1 _5507_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6487_ _6487_/A _6487_/B vssd1 vssd1 vccd1 vccd1 _6487_/X sky130_fd_sc_hd__and2_1
X_8226_ _6353_/A _8225_/X _8223_/Y vssd1 vssd1 vccd1 vccd1 _8226_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_23_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _9650_/CLK sky130_fd_sc_hd__clkbuf_16
X_5438_ _7317_/A vssd1 vssd1 vccd1 vccd1 _7160_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_160_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8157_ _7738_/A _8107_/X _8156_/Y vssd1 vssd1 vccd1 vccd1 _8157_/X sky130_fd_sc_hd__o21ba_1
X_5369_ _5362_/B _5356_/X _5368_/Y _5332_/A _5364_/X vssd1 vssd1 vccd1 vccd1 _5370_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8088_ _9560_/Q vssd1 vssd1 vccd1 vccd1 _8088_/Y sky130_fd_sc_hd__inv_2
X_7108_ _7108_/A _7108_/B vssd1 vssd1 vccd1 vccd1 _7109_/B sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_38_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _9915_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_87_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7039_ _7012_/X _7035_/X _7012_/X _7035_/X vssd1 vssd1 vccd1 vccd1 _7056_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6410_ _9773_/Q _8203_/A _6407_/Y vssd1 vssd1 vccd1 vccd1 _6544_/B sky130_fd_sc_hd__a21oi_2
XFILLER_174_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7390_ _9624_/Q _7408_/B _7467_/A vssd1 vssd1 vccd1 vccd1 _7391_/B sky130_fd_sc_hd__and3_1
XFILLER_174_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6341_ _6341_/A vssd1 vssd1 vccd1 vccd1 _6341_/Y sky130_fd_sc_hd__inv_2
X_6272_ _8031_/A _6143_/X _6268_/X vssd1 vssd1 vccd1 vccd1 _6272_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_170_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9060_ _8028_/Y _8027_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9060_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8011_ _9398_/X _8030_/B vssd1 vssd1 vccd1 vccd1 _8011_/X sky130_fd_sc_hd__and2_1
XFILLER_69_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5223_ _5271_/A vssd1 vssd1 vccd1 vccd1 _5224_/A sky130_fd_sc_hd__clkbuf_2
X_5154_ _9779_/Q _5151_/X input40/X _5152_/X _5153_/X vssd1 vssd1 vccd1 vccd1 _9779_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_130_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5085_ _9803_/Q vssd1 vssd1 vccd1 vccd1 _6318_/A sky130_fd_sc_hd__inv_2
XFILLER_110_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8913_ _8913_/A _8913_/B vssd1 vssd1 vccd1 vccd1 _8913_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9893_ _9893_/CLK _9893_/D vssd1 vssd1 vccd1 vccd1 _9893_/Q sky130_fd_sc_hd__dfxtp_1
X_8844_ _8409_/X _8843_/X _8409_/X _8843_/X vssd1 vssd1 vccd1 vccd1 _8845_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8775_ _8775_/A _8775_/B vssd1 vssd1 vccd1 vccd1 _8781_/A sky130_fd_sc_hd__or2_1
X_5987_ _5987_/A vssd1 vssd1 vccd1 vccd1 _5989_/A sky130_fd_sc_hd__inv_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4938_ _5405_/A vssd1 vssd1 vccd1 vccd1 _4991_/A sky130_fd_sc_hd__clkbuf_4
X_7726_ _7726_/A vssd1 vssd1 vccd1 vccd1 _7726_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7657_ _7657_/A _7657_/B vssd1 vssd1 vccd1 vccd1 _7658_/B sky130_fd_sc_hd__nor2_2
XFILLER_138_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4869_ _9894_/Q _4879_/A _9746_/Q _4880_/A _4867_/X vssd1 vssd1 vccd1 vccd1 _9894_/D
+ sky130_fd_sc_hd__o221a_1
X_6608_ _9464_/X vssd1 vssd1 vccd1 vccd1 _6660_/B sky130_fd_sc_hd__buf_1
XFILLER_192_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7588_ _7588_/A vssd1 vssd1 vccd1 vccd1 _7594_/A sky130_fd_sc_hd__inv_2
X_9327_ _7905_/Y _9778_/Q _9327_/S vssd1 vssd1 vccd1 vccd1 _9327_/X sky130_fd_sc_hd__mux2_1
X_6539_ _6541_/A _6539_/B vssd1 vssd1 vccd1 vccd1 _6539_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9258_ _9257_/X input46/X _9294_/S vssd1 vssd1 vccd1 vccd1 _9258_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8209_ _8231_/B vssd1 vssd1 vccd1 vccd1 _8209_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9189_ _6531_/Y _9794_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9543_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5910_ _5910_/A vssd1 vssd1 vccd1 vccd1 _5915_/A sky130_fd_sc_hd__buf_1
X_6890_ _6890_/A _6890_/B vssd1 vssd1 vccd1 vccd1 _6902_/A sky130_fd_sc_hd__or2_1
X_5841_ _9636_/Q _5832_/X _5039_/X _5833_/X _5840_/X vssd1 vssd1 vccd1 vccd1 _9636_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8560_ _8559_/A _8559_/B _8603_/A vssd1 vssd1 vccd1 vccd1 _8560_/Y sky130_fd_sc_hd__o21ai_1
X_5772_ _5772_/A vssd1 vssd1 vccd1 vccd1 _5772_/X sky130_fd_sc_hd__buf_1
XFILLER_61_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8491_ _8491_/A _8491_/B vssd1 vssd1 vccd1 vccd1 _8526_/A sky130_fd_sc_hd__or2_1
X_7511_ _7503_/A _7503_/B _7503_/X vssd1 vssd1 vccd1 vccd1 _7511_/X sky130_fd_sc_hd__a21bo_1
XFILLER_159_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7442_ _7442_/A _7442_/B vssd1 vssd1 vccd1 vccd1 _7443_/B sky130_fd_sc_hd__nor2_1
XFILLER_147_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7373_ _7294_/X _7372_/Y _7294_/X _7372_/Y vssd1 vssd1 vccd1 vccd1 _7374_/B sky130_fd_sc_hd__a2bb2o_1
X_6324_ _6324_/A _6522_/A vssd1 vssd1 vccd1 vccd1 _6324_/Y sky130_fd_sc_hd__nor2_1
X_9112_ _9596_/Q _5039_/A _9667_/Q vssd1 vssd1 vccd1 vccd1 _9112_/X sky130_fd_sc_hd__mux2_1
X_6255_ _9585_/Q _6169_/A _8027_/A _6245_/A vssd1 vssd1 vccd1 vccd1 _6265_/C sky130_fd_sc_hd__a22o_1
XFILLER_115_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9043_ _7996_/Y _9042_/X _9052_/S vssd1 vssd1 vccd1 vccd1 _9043_/X sky130_fd_sc_hd__mux2_1
X_5206_ _5206_/A vssd1 vssd1 vccd1 vccd1 _5206_/X sky130_fd_sc_hd__clkbuf_2
X_6186_ _9573_/Q _6167_/A _7988_/A _6137_/A vssd1 vssd1 vccd1 vccd1 _6200_/A sky130_fd_sc_hd__a22o_1
X_5137_ _5136_/X _9786_/Q _5130_/X _9213_/X _5132_/X vssd1 vssd1 vccd1 vccd1 _9786_/D
+ sky130_fd_sc_hd__o221a_1
X_5068_ _5061_/X _6317_/A _5067_/Y _5050_/X vssd1 vssd1 vccd1 vccd1 _5069_/B sky130_fd_sc_hd__o22a_1
XFILLER_123_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9876_ _9893_/CLK _9876_/D vssd1 vssd1 vccd1 vccd1 _9876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8827_ _8827_/A vssd1 vssd1 vccd1 vccd1 _8827_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8758_ _8735_/A _8751_/B _8686_/A _8734_/X _8735_/X vssd1 vssd1 vccd1 vccd1 _8826_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7709_ _7877_/A vssd1 vssd1 vccd1 vccd1 _7709_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8689_ _9392_/X vssd1 vssd1 vccd1 vccd1 _8875_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_138_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6040_ _6036_/Y _6039_/X _6036_/Y _6039_/X vssd1 vssd1 vccd1 vccd1 _6040_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7991_ _7991_/A vssd1 vssd1 vccd1 vccd1 _8009_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_39_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9730_ _9879_/CLK _9730_/D vssd1 vssd1 vccd1 vccd1 _9730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6942_ _6941_/A _6941_/B _6941_/X vssd1 vssd1 vccd1 vccd1 _6954_/A sky130_fd_sc_hd__a21boi_1
XFILLER_54_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9661_ _9673_/CLK _9661_/D vssd1 vssd1 vccd1 vccd1 _9661_/Q sky130_fd_sc_hd__dfxtp_1
X_6873_ _9616_/Q _6891_/B _6951_/A vssd1 vssd1 vccd1 vccd1 _6874_/B sky130_fd_sc_hd__and3_1
X_8612_ _8702_/C _8611_/A _8609_/A _8611_/Y vssd1 vssd1 vccd1 vccd1 _8612_/X sky130_fd_sc_hd__a22o_1
X_5824_ _5832_/A vssd1 vssd1 vccd1 vccd1 _5824_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9592_ _9924_/CLK _9592_/D vssd1 vssd1 vccd1 vccd1 _9592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8543_ _8543_/A _8543_/B vssd1 vssd1 vccd1 vccd1 _8626_/C sky130_fd_sc_hd__nor2_4
XFILLER_148_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5755_ _9680_/Q _9663_/Q _5716_/Y _5754_/X vssd1 vssd1 vccd1 vccd1 _5755_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_10_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8474_ _9378_/X vssd1 vssd1 vccd1 vccd1 _8584_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_175_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5686_ _6576_/A _5681_/X _9104_/X _5684_/X _5682_/X vssd1 vssd1 vccd1 vccd1 _9677_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7425_ _7378_/X _7423_/X _7378_/X _7423_/X vssd1 vssd1 vccd1 vccd1 _7425_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_190_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7356_ _7332_/X _7353_/X _7332_/X _7353_/X vssd1 vssd1 vccd1 vccd1 _7356_/X sky130_fd_sc_hd__a2bb2o_1
X_6307_ _9844_/Q _6486_/A _4976_/X _6487_/A vssd1 vssd1 vccd1 vccd1 _6307_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7287_ _7276_/A _7276_/B _7276_/X vssd1 vssd1 vccd1 vccd1 _7288_/B sky130_fd_sc_hd__a21bo_1
X_6238_ _8017_/A _6193_/X _6244_/A _6234_/X vssd1 vssd1 vccd1 vccd1 _6238_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9026_ _7965_/Y _9601_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9026_/X sky130_fd_sc_hd__mux2_1
X_6169_ _6169_/A vssd1 vssd1 vccd1 vccd1 _6170_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9928_ _9928_/CLK _9928_/D vssd1 vssd1 vccd1 vccd1 _9928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9859_ _9930_/CLK _9859_/D vssd1 vssd1 vccd1 vccd1 _9859_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5540_ _9394_/X _5481_/X _5482_/X _5539_/X vssd1 vssd1 vccd1 vccd1 _5566_/B sky130_fd_sc_hd__o22a_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5471_ _5471_/A vssd1 vssd1 vccd1 vccd1 _5471_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7210_ _7210_/A _7210_/B _7210_/C vssd1 vssd1 vccd1 vccd1 _7506_/A sky130_fd_sc_hd__and3_1
XFILLER_144_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8190_ _9847_/Q _6360_/Y _8183_/Y _8189_/X vssd1 vssd1 vccd1 vccd1 _8191_/B sky130_fd_sc_hd__o22a_1
XFILLER_125_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7141_ _7386_/A vssd1 vssd1 vccd1 vccd1 _7394_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7072_ _7072_/A _7072_/B vssd1 vssd1 vccd1 vccd1 _7073_/B sky130_fd_sc_hd__or2_1
X_6023_ _9641_/Q vssd1 vssd1 vccd1 vccd1 _6023_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7974_ _7974_/A _7981_/B vssd1 vssd1 vccd1 vccd1 _7974_/X sky130_fd_sc_hd__or2_1
XFILLER_82_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9713_ _9828_/CLK _9713_/D vssd1 vssd1 vccd1 vccd1 _9713_/Q sky130_fd_sc_hd__dfxtp_1
X_6925_ _6925_/A _6925_/B vssd1 vssd1 vccd1 vccd1 _6926_/B sky130_fd_sc_hd__nor2_1
XPHY_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9644_ _9650_/CLK _9644_/D vssd1 vssd1 vccd1 vccd1 _9644_/Q sky130_fd_sc_hd__dfxtp_1
X_6856_ _6777_/X _6855_/Y _6777_/X _6855_/Y vssd1 vssd1 vccd1 vccd1 _6857_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5807_ _5744_/A _5806_/Y _5744_/A _5806_/Y vssd1 vssd1 vccd1 vccd1 _5808_/A sky130_fd_sc_hd__a2bb2o_1
X_9575_ _9578_/CLK _9575_/D vssd1 vssd1 vccd1 vccd1 _9575_/Q sky130_fd_sc_hd__dfxtp_1
X_6787_ _6787_/A _6855_/B vssd1 vssd1 vccd1 vccd1 _6787_/Y sky130_fd_sc_hd__nor2_1
XFILLER_195_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8526_ _8526_/A _8526_/B vssd1 vssd1 vccd1 vccd1 _8559_/A sky130_fd_sc_hd__nor2_2
X_5738_ _9655_/Q vssd1 vssd1 vccd1 vccd1 _5738_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8457_ _8457_/A _8457_/B vssd1 vssd1 vccd1 vccd1 _8458_/A sky130_fd_sc_hd__or2_1
XFILLER_135_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5669_ _9669_/Q vssd1 vssd1 vccd1 vccd1 _6571_/A sky130_fd_sc_hd__buf_2
XFILLER_190_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8388_ _9691_/Q vssd1 vssd1 vccd1 vccd1 _8389_/A sky130_fd_sc_hd__inv_2
X_7408_ _9626_/Q _7408_/B _7419_/A vssd1 vssd1 vccd1 vccd1 _7409_/A sky130_fd_sc_hd__and3_1
XFILLER_150_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7339_ _7330_/A _7336_/Y _7337_/X _7338_/X vssd1 vssd1 vccd1 vccd1 _7352_/B sky130_fd_sc_hd__o22ai_2
XFILLER_131_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9009_ _9564_/Q _9522_/Q _9013_/S vssd1 vssd1 vccd1 vccd1 _9009_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4971_ _4960_/X _9445_/S _4965_/A _4970_/X _4955_/X vssd1 vssd1 vccd1 vccd1 _9847_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7690_ _8134_/A _8184_/B _7901_/A _9777_/Q _7689_/X vssd1 vssd1 vccd1 vccd1 _7705_/A
+ sky130_fd_sc_hd__o221a_1
X_6710_ _9094_/X vssd1 vssd1 vccd1 vccd1 _6756_/B sky130_fd_sc_hd__inv_2
X_6641_ _9463_/X vssd1 vssd1 vccd1 vccd1 _6691_/B sky130_fd_sc_hd__inv_2
XFILLER_177_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9360_ _7613_/X _7581_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9360_/X sky130_fd_sc_hd__mux2_2
XFILLER_192_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8311_ _7696_/X _9540_/Q _7755_/X _9539_/Q vssd1 vssd1 vccd1 vccd1 _8311_/X sky130_fd_sc_hd__o22a_1
X_6572_ _6867_/C vssd1 vssd1 vccd1 vccd1 _6890_/A sky130_fd_sc_hd__clkbuf_4
X_5523_ _5617_/A _5617_/B vssd1 vssd1 vccd1 vccd1 _5616_/A sky130_fd_sc_hd__nand2_1
XFILLER_145_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9291_ _7859_/Y _9768_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9291_/X sky130_fd_sc_hd__mux2_1
X_8242_ _6337_/A _8240_/B _8240_/X vssd1 vssd1 vccd1 vccd1 _8242_/X sky130_fd_sc_hd__a21bo_1
X_5454_ _9337_/X _9336_/X _5428_/X _5453_/X vssd1 vssd1 vccd1 vccd1 _5454_/X sky130_fd_sc_hd__o22a_1
X_8173_ _8174_/A _8174_/B _8172_/Y vssd1 vssd1 vccd1 vccd1 _8175_/A sky130_fd_sc_hd__a21oi_1
XFILLER_172_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5385_ _9721_/Q _5385_/B vssd1 vssd1 vccd1 vccd1 _5385_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7124_ _5764_/Y _7121_/X _5764_/Y _7121_/X vssd1 vssd1 vccd1 vccd1 _7124_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7055_ _7055_/A vssd1 vssd1 vccd1 vccd1 _7055_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6006_ _7941_/A _9638_/Q _5998_/B _6001_/X vssd1 vssd1 vccd1 vccd1 _6006_/X sky130_fd_sc_hd__o22a_1
XFILLER_55_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7957_ _7957_/A _9013_/S vssd1 vssd1 vccd1 vccd1 _7957_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7888_ _7680_/A _7883_/Y _7860_/X _7892_/B vssd1 vssd1 vccd1 vccd1 _7888_/X sky130_fd_sc_hd__o211a_1
X_6908_ _6861_/X _6906_/X _6861_/X _6906_/X vssd1 vssd1 vccd1 vccd1 _6908_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9627_ _9634_/CLK _9627_/D vssd1 vssd1 vccd1 vccd1 _9627_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6839_ _6815_/X _6836_/X _6815_/X _6836_/X vssd1 vssd1 vccd1 vccd1 _6839_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_210_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9558_ _9928_/CLK _9558_/D vssd1 vssd1 vccd1 vccd1 _9558_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8509_ _8576_/C _8472_/X _8473_/X _8476_/X vssd1 vssd1 vccd1 vccd1 _8531_/B sky130_fd_sc_hd__o22ai_4
X_9489_ _9488_/X _6969_/A _9507_/S vssd1 vssd1 vccd1 vccd1 _9489_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_4_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _9833_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5170_ _9772_/Q vssd1 vssd1 vccd1 vccd1 _6347_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_142_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput4 io_wb_adr_i[10] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_1
X_8860_ _8859_/A _8859_/B _8859_/X vssd1 vssd1 vccd1 vccd1 _8927_/A sky130_fd_sc_hd__a21bo_1
XFILLER_64_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8791_ _8749_/X _8790_/X _8749_/X _8790_/X vssd1 vssd1 vccd1 vccd1 _8792_/A sky130_fd_sc_hd__a2bb2o_1
X_7811_ _7769_/A _7810_/B _7785_/X _7814_/B vssd1 vssd1 vccd1 vccd1 _7811_/X sky130_fd_sc_hd__o211a_1
XFILLER_91_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7742_ _7844_/A vssd1 vssd1 vccd1 vccd1 _7743_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4954_ _9115_/X _4951_/X _9852_/Q _4952_/X _4947_/X vssd1 vssd1 vccd1 vccd1 _9852_/D
+ sky130_fd_sc_hd__o221a_1
X_7673_ _7673_/A _7673_/B vssd1 vssd1 vccd1 vccd1 _7854_/A sky130_fd_sc_hd__or2_1
X_9412_ _9411_/X _7490_/A _9506_/S vssd1 vssd1 vccd1 vccd1 _9412_/X sky130_fd_sc_hd__mux2_1
X_4885_ _9737_/Q _4879_/X _9885_/Q _4880_/X _4881_/X vssd1 vssd1 vccd1 vccd1 _9885_/D
+ sky130_fd_sc_hd__a221o_1
X_6624_ _9461_/X vssd1 vssd1 vccd1 vccd1 _6969_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_177_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6555_ _9672_/Q _6565_/A vssd1 vssd1 vccd1 vccd1 _6556_/B sky130_fd_sc_hd__or2_1
X_9343_ _7629_/X _7589_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9343_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5506_ _9380_/X _5505_/X _9380_/X _5505_/X vssd1 vssd1 vccd1 vccd1 _5612_/A sky130_fd_sc_hd__a2bb2oi_1
X_9274_ _9273_/X input19/X _9282_/S vssd1 vssd1 vccd1 vccd1 _9274_/X sky130_fd_sc_hd__mux2_1
X_6486_ _6486_/A _6486_/B vssd1 vssd1 vccd1 vccd1 _6486_/X sky130_fd_sc_hd__or2_1
XFILLER_118_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8225_ _8225_/A _8227_/B vssd1 vssd1 vccd1 vccd1 _8225_/X sky130_fd_sc_hd__or2_1
XFILLER_133_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5437_ _7314_/A vssd1 vssd1 vccd1 vccd1 _7317_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8156_ _7723_/A _8108_/X _8155_/X vssd1 vssd1 vccd1 vccd1 _8156_/Y sky130_fd_sc_hd__o21ai_1
X_5368_ _9725_/Q _5368_/B vssd1 vssd1 vccd1 vccd1 _5368_/Y sky130_fd_sc_hd__nor2_1
X_8087_ _8089_/B vssd1 vssd1 vccd1 vccd1 _8087_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7107_ _7107_/A _7107_/B vssd1 vssd1 vccd1 vccd1 _7108_/B sky130_fd_sc_hd__or2_1
X_5299_ _9736_/Q _5299_/B vssd1 vssd1 vccd1 vccd1 _5299_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7038_ _6968_/X _7037_/X _6968_/X _7037_/X vssd1 vssd1 vccd1 vccd1 _7038_/Y sky130_fd_sc_hd__a2bb2oi_2
XFILLER_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8989_ _8988_/X _7490_/A _9506_/S vssd1 vssd1 vccd1 vccd1 _8989_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6340_ _9788_/Q vssd1 vssd1 vccd1 vccd1 _6340_/Y sky130_fd_sc_hd__inv_2
X_6271_ _9588_/Q _6170_/A _8033_/A _6141_/A vssd1 vssd1 vccd1 vccd1 _6271_/X sky130_fd_sc_hd__a22o_1
XFILLER_115_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5222_ _5222_/A _5919_/A vssd1 vssd1 vccd1 vccd1 _5271_/A sky130_fd_sc_hd__or2_2
X_8010_ _8010_/A _8010_/B vssd1 vssd1 vccd1 vccd1 _8010_/Y sky130_fd_sc_hd__nor2_1
X_5153_ _5165_/A vssd1 vssd1 vccd1 vccd1 _5153_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5084_ _5136_/A vssd1 vssd1 vccd1 vccd1 _5084_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8912_ _8935_/A _9422_/X _8820_/X vssd1 vssd1 vccd1 vccd1 _8913_/B sky130_fd_sc_hd__or3b_1
X_9892_ _9893_/CLK _9892_/D vssd1 vssd1 vccd1 vccd1 _9892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8843_ _8381_/A _6593_/A _8381_/Y vssd1 vssd1 vccd1 vccd1 _8843_/X sky130_fd_sc_hd__a21o_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8774_ _8774_/A vssd1 vssd1 vccd1 vccd1 _8775_/B sky130_fd_sc_hd__inv_2
X_5986_ _7935_/A _9637_/Q _9850_/Q _5985_/Y vssd1 vssd1 vccd1 vccd1 _5987_/A sky130_fd_sc_hd__o22a_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7725_ _7814_/A vssd1 vssd1 vccd1 vccd1 _7726_/A sky130_fd_sc_hd__clkbuf_2
X_4937_ _9125_/X _4934_/X _9862_/Q _4935_/X _4923_/X vssd1 vssd1 vccd1 vccd1 _9862_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7656_ _9899_/Q _7777_/A vssd1 vssd1 vccd1 vccd1 _7657_/B sky130_fd_sc_hd__or2_2
XFILLER_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4868_ _9895_/Q _4865_/X _9747_/Q _4866_/X _4867_/X vssd1 vssd1 vccd1 vccd1 _9895_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_192_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6607_ _6706_/A vssd1 vssd1 vccd1 vccd1 _6969_/A sky130_fd_sc_hd__buf_2
XFILLER_20_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9326_ _9325_/X input37/X _9334_/S vssd1 vssd1 vccd1 vccd1 _9326_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4799_ _4799_/A vssd1 vssd1 vccd1 vccd1 _4799_/X sky130_fd_sc_hd__buf_2
X_7587_ _7587_/A vssd1 vssd1 vccd1 vccd1 _7595_/A sky130_fd_sc_hd__inv_2
XFILLER_146_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6538_ _6541_/A _6538_/B vssd1 vssd1 vccd1 vccd1 _6538_/Y sky130_fd_sc_hd__nor2_1
XFILLER_161_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6469_ _9755_/Q vssd1 vssd1 vccd1 vccd1 _6469_/Y sky130_fd_sc_hd__inv_2
X_9257_ _9256_/X _7811_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9257_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8208_ _8204_/A _8204_/B _8205_/B vssd1 vssd1 vccd1 vccd1 _8208_/Y sky130_fd_sc_hd__o21ai_1
X_9188_ _6529_/Y _9793_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9542_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8139_ _7803_/A _8121_/X _7707_/A _8120_/X _8138_/X vssd1 vssd1 vccd1 vccd1 _8139_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_121_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _9828_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_179_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5840_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5840_/X sky130_fd_sc_hd__buf_2
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5771_ _5754_/X _5770_/X _5754_/X _5770_/X vssd1 vssd1 vccd1 vccd1 _7120_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_194_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8490_ _8491_/B vssd1 vssd1 vccd1 vccd1 _8490_/Y sky130_fd_sc_hd__inv_2
X_7510_ _7506_/X _7507_/X _7506_/X _7507_/X vssd1 vssd1 vccd1 vccd1 _7514_/A sky130_fd_sc_hd__a2bb2o_1
X_7441_ _7415_/A _7421_/A _7415_/Y vssd1 vssd1 vccd1 vccd1 _7441_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_37_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _9578_/CLK sky130_fd_sc_hd__clkbuf_16
Xinput40 io_wb_dat_i[31] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7372_ _7372_/A _7372_/B vssd1 vssd1 vccd1 vccd1 _7372_/Y sky130_fd_sc_hd__nor2_1
X_6323_ _6542_/A vssd1 vssd1 vccd1 vccd1 _6522_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9111_ _9595_/Q _5041_/A _9667_/Q vssd1 vssd1 vccd1 vccd1 _9111_/X sky130_fd_sc_hd__mux2_1
X_6254_ _9585_/Q vssd1 vssd1 vccd1 vccd1 _8027_/A sky130_fd_sc_hd__inv_2
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9042_ _7997_/Y _9607_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9042_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5205_ _5205_/A vssd1 vssd1 vccd1 vccd1 _5205_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6185_ _9573_/Q vssd1 vssd1 vccd1 vccd1 _7988_/A sky130_fd_sc_hd__inv_2
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5136_ _5136_/A vssd1 vssd1 vccd1 vccd1 _5136_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5067_ _9839_/Q vssd1 vssd1 vccd1 vccd1 _5067_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9875_ _9893_/CLK _9875_/D vssd1 vssd1 vccd1 vccd1 _9875_/Q sky130_fd_sc_hd__dfxtp_1
X_8826_ _8826_/A _8757_/X vssd1 vssd1 vccd1 vccd1 _8827_/A sky130_fd_sc_hd__or2b_1
X_8757_ _5858_/X _8754_/Y _8755_/X _8756_/Y vssd1 vssd1 vccd1 vccd1 _8757_/X sky130_fd_sc_hd__a31o_1
X_5969_ _9518_/D vssd1 vssd1 vccd1 vccd1 _5969_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7708_ _9921_/Q vssd1 vssd1 vccd1 vccd1 _7877_/A sky130_fd_sc_hd__inv_2
X_8688_ _8751_/B vssd1 vssd1 vccd1 vccd1 _8958_/B sky130_fd_sc_hd__buf_1
XFILLER_193_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7639_ _7639_/A _7640_/B vssd1 vssd1 vccd1 vccd1 _7639_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9309_ _9308_/X _7884_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9309_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7990_ _7990_/A _8003_/B vssd1 vssd1 vccd1 vccd1 _7990_/X sky130_fd_sc_hd__or2_1
XFILLER_93_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6941_ _6941_/A _6941_/B vssd1 vssd1 vccd1 vccd1 _6941_/X sky130_fd_sc_hd__or2_1
XFILLER_207_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9660_ _9673_/CLK _9660_/D vssd1 vssd1 vccd1 vccd1 _9660_/Q sky130_fd_sc_hd__dfxtp_1
X_6872_ _6872_/A _6872_/B vssd1 vssd1 vccd1 vccd1 _6951_/A sky130_fd_sc_hd__or2_2
XFILLER_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8611_ _8611_/A vssd1 vssd1 vccd1 vccd1 _8611_/Y sky130_fd_sc_hd__inv_2
X_9591_ _9924_/CLK _9591_/D vssd1 vssd1 vccd1 vccd1 _9591_/Q sky130_fd_sc_hd__dfxtp_1
X_5823_ _9648_/Q _5818_/X input20/X _5819_/X _5822_/X vssd1 vssd1 vccd1 vccd1 _9648_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_62_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8542_ _8540_/X _8541_/X _8540_/X _8541_/X vssd1 vssd1 vccd1 vccd1 _8542_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_194_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5754_ _5717_/Y _5718_/Y _5719_/X _5753_/X vssd1 vssd1 vccd1 vccd1 _5754_/X sky130_fd_sc_hd__o22a_1
X_8473_ _8576_/C _8472_/X _8576_/C _8472_/X vssd1 vssd1 vccd1 vccd1 _8473_/X sky130_fd_sc_hd__a2bb2o_2
X_5685_ _6577_/A _5681_/X _9105_/X _5684_/X _5682_/X vssd1 vssd1 vccd1 vccd1 _9678_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7424_ _7260_/A _7260_/B _7427_/B vssd1 vssd1 vccd1 vccd1 _7424_/X sky130_fd_sc_hd__a21o_1
X_7355_ _7307_/X _7354_/X _7307_/X _7354_/X vssd1 vssd1 vccd1 vccd1 _7355_/X sky130_fd_sc_hd__a2bb2o_1
X_6306_ _9781_/Q vssd1 vssd1 vccd1 vccd1 _6486_/A sky130_fd_sc_hd__inv_2
XFILLER_103_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7286_ _7286_/A _7267_/X vssd1 vssd1 vccd1 vccd1 _7288_/A sky130_fd_sc_hd__or2b_1
XFILLER_131_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6237_ _9582_/Q _6169_/A _8019_/A _6139_/A vssd1 vssd1 vccd1 vccd1 _6244_/B sky130_fd_sc_hd__a22o_1
X_9025_ _9024_/X _9754_/Q _9481_/S vssd1 vssd1 vccd1 vccd1 _9025_/X sky130_fd_sc_hd__mux2_2
X_6168_ _6168_/A vssd1 vssd1 vccd1 vccd1 _6169_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_134_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5119_ _5128_/A _6500_/A _5118_/Y _5097_/A vssd1 vssd1 vccd1 vccd1 _5120_/B sky130_fd_sc_hd__o22a_1
XFILLER_57_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6099_ _6095_/X _6098_/X _6095_/X _6098_/X vssd1 vssd1 vccd1 vccd1 _6099_/X sky130_fd_sc_hd__o2bb2a_1
X_9927_ _9928_/CLK _9927_/D vssd1 vssd1 vccd1 vccd1 _9927_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_150_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9858_ _9858_/CLK _9858_/D vssd1 vssd1 vccd1 vccd1 _9858_/Q sky130_fd_sc_hd__dfxtp_1
X_8809_ _8804_/X _8808_/X _8804_/X _8808_/X vssd1 vssd1 vccd1 vccd1 _8812_/A sky130_fd_sc_hd__a2bb2oi_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9789_ _9929_/CLK _9789_/D vssd1 vssd1 vccd1 vccd1 _9789_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5470_ _9420_/X _5469_/X _9420_/X _5469_/X vssd1 vssd1 vccd1 vccd1 _5555_/A sky130_fd_sc_hd__a2bb2oi_1
XFILLER_172_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7140_ _9624_/Q vssd1 vssd1 vccd1 vccd1 _7386_/A sky130_fd_sc_hd__inv_2
X_7071_ _7071_/A _7071_/B vssd1 vssd1 vccd1 vccd1 _7072_/B sky130_fd_sc_hd__or2_1
XFILLER_100_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6022_ _6018_/A _6021_/X _6018_/A _6021_/X vssd1 vssd1 vccd1 vccd1 _6022_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_100_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7973_ _7973_/A _7993_/B vssd1 vssd1 vccd1 vccd1 _7973_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9712_ _9828_/CLK _9712_/D vssd1 vssd1 vccd1 vccd1 _9712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6924_ _6898_/A _6904_/A _6898_/Y vssd1 vssd1 vccd1 vccd1 _6924_/X sky130_fd_sc_hd__a21o_1
XPHY_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9643_ _9650_/CLK _9643_/D vssd1 vssd1 vccd1 vccd1 _9643_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6855_ _6855_/A _6855_/B vssd1 vssd1 vccd1 vccd1 _6855_/Y sky130_fd_sc_hd__nor2_2
XFILLER_210_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5806_ _9670_/Q _9653_/Q _5741_/Y vssd1 vssd1 vccd1 vccd1 _5806_/Y sky130_fd_sc_hd__a21oi_1
X_9574_ _9909_/CLK _9574_/D vssd1 vssd1 vccd1 vccd1 _9574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6786_ _6786_/A _6786_/B vssd1 vssd1 vccd1 vccd1 _6855_/B sky130_fd_sc_hd__nor2_2
XFILLER_210_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8525_ _8525_/A vssd1 vssd1 vccd1 vccd1 _8526_/B sky130_fd_sc_hd__inv_2
XFILLER_148_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5737_ _9672_/Q vssd1 vssd1 vccd1 vccd1 _6564_/A sky130_fd_sc_hd__inv_2
X_8456_ _8455_/A _8455_/B _8455_/Y vssd1 vssd1 vccd1 vccd1 _8457_/B sky130_fd_sc_hd__a21o_1
XFILLER_148_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5668_ _9686_/Q _5658_/X _6569_/A _5662_/X _5660_/X vssd1 vssd1 vccd1 vccd1 _9686_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_108_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7407_ _7407_/A _7407_/B vssd1 vssd1 vccd1 vccd1 _7419_/A sky130_fd_sc_hd__or2_1
X_5599_ _5599_/A vssd1 vssd1 vccd1 vccd1 _5599_/Y sky130_fd_sc_hd__inv_2
X_8387_ _9692_/Q _6582_/X _9692_/Q _6582_/X vssd1 vssd1 vccd1 vccd1 _8387_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_190_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7338_ _7323_/X _7324_/X _7323_/X _7324_/X vssd1 vssd1 vccd1 vccd1 _7338_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_145_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7269_ _7324_/A _9470_/X vssd1 vssd1 vccd1 vccd1 _7269_/X sky130_fd_sc_hd__or2_1
X_9008_ _9007_/X _9749_/Q _9481_/S vssd1 vssd1 vccd1 vccd1 _9008_/X sky130_fd_sc_hd__mux2_4
XFILLER_77_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_20 _9930_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4970_ _4969_/A _4969_/B _4968_/Y _5026_/A _4969_/Y vssd1 vssd1 vccd1 vccd1 _4970_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_91_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6640_ _6678_/A _9462_/X vssd1 vssd1 vccd1 vccd1 _6647_/C sky130_fd_sc_hd__nor2_1
X_6571_ _6571_/A vssd1 vssd1 vccd1 vccd1 _6571_/Y sky130_fd_sc_hd__inv_2
X_5522_ _9446_/X _5509_/X _9446_/X _5509_/X vssd1 vssd1 vccd1 vccd1 _5617_/B sky130_fd_sc_hd__a2bb2oi_1
X_8310_ _7769_/Y _9537_/Q _7726_/X _9538_/Q vssd1 vssd1 vccd1 vccd1 _8310_/X sky130_fd_sc_hd__o22a_1
XFILLER_185_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9290_ _9289_/X input25/X _9294_/S vssd1 vssd1 vccd1 vccd1 _9290_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8241_ _5198_/X _8240_/X _8232_/B vssd1 vssd1 vccd1 vccd1 _8241_/X sky130_fd_sc_hd__a21bo_1
XFILLER_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5453_ _9343_/X _9341_/X _5431_/Y _5503_/A vssd1 vssd1 vccd1 vccd1 _5453_/X sky130_fd_sc_hd__o22a_1
X_8172_ _4770_/X _8091_/X _8171_/X vssd1 vssd1 vccd1 vccd1 _8172_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_160_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5384_ _5384_/A vssd1 vssd1 vccd1 vccd1 _5385_/B sky130_fd_sc_hd__inv_2
X_7123_ _7120_/A _7120_/B _7121_/B vssd1 vssd1 vccd1 vccd1 _7123_/X sky130_fd_sc_hd__a21bo_1
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7054_ _7054_/A _7054_/B vssd1 vssd1 vccd1 vccd1 _7055_/A sky130_fd_sc_hd__or2_1
X_6005_ _7947_/A _9639_/Q _9852_/Q _6004_/Y vssd1 vssd1 vccd1 vccd1 _6008_/A sky130_fd_sc_hd__a22o_1
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7956_ _9502_/X _7956_/B vssd1 vssd1 vccd1 vccd1 _7956_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7887_ _7887_/A _7887_/B vssd1 vssd1 vccd1 vccd1 _7892_/B sky130_fd_sc_hd__or2_2
X_6907_ _6743_/A _6743_/B _6910_/B vssd1 vssd1 vccd1 vccd1 _6907_/X sky130_fd_sc_hd__a21o_1
XFILLER_35_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9626_ _9858_/CLK _9626_/D vssd1 vssd1 vccd1 vccd1 _9626_/Q sky130_fd_sc_hd__dfxtp_2
X_6838_ _6790_/X _6837_/X _6790_/X _6837_/X vssd1 vssd1 vccd1 vccd1 _6838_/X sky130_fd_sc_hd__a2bb2o_1
X_9557_ _9924_/CLK _9557_/D vssd1 vssd1 vccd1 vccd1 _9557_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_8508_ _8508_/A vssd1 vssd1 vccd1 vccd1 _8510_/A sky130_fd_sc_hd__inv_2
XFILLER_136_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6769_ _6769_/A _6750_/X vssd1 vssd1 vccd1 vccd1 _6771_/A sky130_fd_sc_hd__or2b_1
XFILLER_148_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9488_ _9487_/X _7494_/A _9506_/S vssd1 vssd1 vccd1 vccd1 _9488_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8439_ _8472_/C _8438_/B _8460_/A vssd1 vssd1 vccd1 vccd1 _8441_/B sky130_fd_sc_hd__o21ai_2
XFILLER_136_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput5 io_wb_adr_i[11] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_1
X_7810_ _7810_/A _7810_/B vssd1 vssd1 vccd1 vccd1 _7814_/B sky130_fd_sc_hd__nand2_2
X_8790_ _8763_/X _8789_/X _8763_/X _8789_/X vssd1 vssd1 vccd1 vccd1 _8790_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7741_ _9913_/Q vssd1 vssd1 vccd1 vccd1 _7844_/A sky130_fd_sc_hd__inv_2
X_4953_ _9116_/X _4951_/X _9853_/Q _4952_/X _4947_/X vssd1 vssd1 vccd1 vccd1 _9853_/D
+ sky130_fd_sc_hd__o221a_1
X_7672_ _9915_/Q _7846_/A vssd1 vssd1 vccd1 vccd1 _7673_/B sky130_fd_sc_hd__or2_2
X_6623_ _9617_/Q _6610_/Y _5890_/X _6612_/Y _6622_/Y vssd1 vssd1 vccd1 vccd1 _6623_/X
+ sky130_fd_sc_hd__a41o_1
X_9411_ _9410_/X _8955_/A _9505_/S vssd1 vssd1 vccd1 vccd1 _9411_/X sky130_fd_sc_hd__mux2_1
X_4884_ _9738_/Q _4879_/X _9886_/Q _4880_/X _4881_/X vssd1 vssd1 vccd1 vccd1 _9886_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6554_ _6567_/A _6554_/B vssd1 vssd1 vccd1 vccd1 _6565_/A sky130_fd_sc_hd__or2_1
X_9342_ _7057_/A _7608_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9342_/X sky130_fd_sc_hd__mux2_1
X_6485_ _9780_/Q _6324_/A _6486_/A _6486_/B vssd1 vssd1 vccd1 vccd1 _6485_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_118_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9273_ _9272_/X _7828_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9273_/X sky130_fd_sc_hd__mux2_1
X_5505_ _5503_/Y _5504_/Y _5503_/Y _5504_/Y vssd1 vssd1 vccd1 vccd1 _5505_/X sky130_fd_sc_hd__a2bb2o_4
X_8224_ _6352_/Y _8223_/Y _8221_/X vssd1 vssd1 vccd1 vccd1 _8224_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5436_ _9619_/Q vssd1 vssd1 vccd1 vccd1 _7314_/A sky130_fd_sc_hd__inv_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8155_ _7723_/A _8108_/X _8154_/Y vssd1 vssd1 vccd1 vccd1 _8155_/X sky130_fd_sc_hd__a21bo_1
XFILLER_99_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5367_ _5367_/A vssd1 vssd1 vccd1 vccd1 _5368_/B sky130_fd_sc_hd__inv_2
X_8086_ _9558_/Q _8093_/A vssd1 vssd1 vccd1 vccd1 _8089_/B sky130_fd_sc_hd__or2_1
XFILLER_141_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5298_ _5298_/A vssd1 vssd1 vccd1 vccd1 _5299_/B sky130_fd_sc_hd__inv_2
X_7106_ _7487_/C vssd1 vssd1 vccd1 vccd1 _7518_/A sky130_fd_sc_hd__buf_2
X_7037_ _7009_/X _7036_/Y _7009_/X _7036_/Y vssd1 vssd1 vccd1 vccd1 _7037_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8988_ _8987_/X _8955_/A _9505_/S vssd1 vssd1 vccd1 vccd1 _8988_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7939_ _8576_/A vssd1 vssd1 vccd1 vccd1 _8865_/A sky130_fd_sc_hd__buf_2
XFILLER_15_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9609_ _9761_/CLK _9609_/D vssd1 vssd1 vccd1 vccd1 _9609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6270_ _9588_/Q vssd1 vssd1 vccd1 vccd1 _8033_/A sky130_fd_sc_hd__inv_2
XFILLER_142_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5221_ _9335_/X vssd1 vssd1 vccd1 vccd1 _5919_/A sky130_fd_sc_hd__inv_2
X_5152_ _5179_/A vssd1 vssd1 vccd1 vccd1 _5152_/X sky130_fd_sc_hd__buf_2
XFILLER_123_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5083_ _5092_/A _5083_/B vssd1 vssd1 vccd1 vccd1 _9804_/D sky130_fd_sc_hd__nor2_1
XFILLER_84_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8911_ _9629_/Q _8908_/Y _5860_/X _8909_/Y _8910_/X vssd1 vssd1 vccd1 vccd1 _8913_/A
+ sky130_fd_sc_hd__a41o_1
X_9891_ _9893_/CLK _9891_/D vssd1 vssd1 vccd1 vccd1 _9891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8842_ _8841_/A _8841_/B _8887_/A vssd1 vssd1 vccd1 vccd1 _8842_/X sky130_fd_sc_hd__a21bo_1
XFILLER_112_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8773_ _8773_/A _8773_/B _8773_/C _8773_/D vssd1 vssd1 vccd1 vccd1 _8774_/A sky130_fd_sc_hd__or4_4
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7724_ _9906_/Q vssd1 vssd1 vccd1 vccd1 _7814_/A sky130_fd_sc_hd__inv_2
X_5985_ _9637_/Q vssd1 vssd1 vccd1 vccd1 _5985_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4936_ _9126_/X _4934_/X _9863_/Q _4935_/X _4923_/X vssd1 vssd1 vccd1 vccd1 _9863_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_193_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7655_ _7749_/A _7776_/A vssd1 vssd1 vccd1 vccd1 _7777_/A sky130_fd_sc_hd__or2_1
X_4867_ _4923_/A vssd1 vssd1 vccd1 vccd1 _4867_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_177_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6606_ _6868_/A vssd1 vssd1 vccd1 vccd1 _6706_/A sky130_fd_sc_hd__buf_1
XFILLER_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7586_ _7586_/A vssd1 vssd1 vccd1 vccd1 _7596_/A sky130_fd_sc_hd__inv_2
X_9325_ _9324_/X _7904_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9325_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4798_ _4798_/A vssd1 vssd1 vccd1 vccd1 _4798_/X sky130_fd_sc_hd__clkbuf_2
X_6537_ _6541_/A _6537_/B vssd1 vssd1 vccd1 vccd1 _6537_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6468_ _8236_/A _6372_/B _6467_/Y vssd1 vssd1 vccd1 vccd1 _6520_/B sky130_fd_sc_hd__a21oi_2
X_9256_ _9756_/Q _9255_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9256_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6399_ _6550_/B vssd1 vssd1 vccd1 vccd1 _6399_/Y sky130_fd_sc_hd__inv_2
X_8207_ _8205_/A _8205_/B _8205_/X vssd1 vssd1 vccd1 vccd1 _8207_/X sky130_fd_sc_hd__a21bo_1
XFILLER_133_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9187_ _6528_/Y _9792_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9541_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5419_ _9353_/X _9351_/X _9353_/X _9351_/X vssd1 vssd1 vccd1 vccd1 _5419_/X sky130_fd_sc_hd__a2bb2o_2
X_8138_ _8123_/Y _8137_/Y _7801_/A _8121_/X vssd1 vssd1 vccd1 vccd1 _8138_/X sky130_fd_sc_hd__a22o_1
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8069_ _9541_/Q _8069_/B vssd1 vssd1 vccd1 vccd1 _8070_/B sky130_fd_sc_hd__or2_1
XFILLER_87_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _9916_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_203_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5770_ _6596_/A _9663_/Q _5716_/Y vssd1 vssd1 vccd1 vccd1 _5770_/X sky130_fd_sc_hd__a21o_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7440_ _7376_/B _7439_/Y _7376_/B _7439_/Y vssd1 vssd1 vccd1 vccd1 _7440_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput30 io_wb_dat_i[22] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9110_ _6112_/X _6114_/X _9896_/Q vssd1 vssd1 vccd1 vccd1 _9110_/X sky130_fd_sc_hd__mux2_1
Xinput41 io_wb_dat_i[3] vssd1 vssd1 vccd1 vccd1 _5035_/A sky130_fd_sc_hd__buf_6
X_7371_ _7307_/X _7354_/X _7355_/X _7370_/X vssd1 vssd1 vccd1 vccd1 _7374_/A sky130_fd_sc_hd__o22a_1
XFILLER_162_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6322_ _9748_/Q vssd1 vssd1 vccd1 vccd1 _6324_/A sky130_fd_sc_hd__inv_2
XFILLER_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6253_ _6265_/B _6252_/X _6265_/B _6252_/X vssd1 vssd1 vccd1 vccd1 _6253_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_88_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9041_ _7994_/X _9040_/X _9053_/S vssd1 vssd1 vccd1 vccd1 _9041_/X sky130_fd_sc_hd__mux2_2
X_5204_ _9756_/Q vssd1 vssd1 vccd1 vccd1 _6341_/A sky130_fd_sc_hd__buf_2
XFILLER_88_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6184_ _6187_/B _6183_/Y _6187_/B _6183_/Y vssd1 vssd1 vccd1 vccd1 _6184_/X sky130_fd_sc_hd__a2bb2o_1
X_5135_ _5128_/X _9787_/Q _5130_/X _9214_/X _5132_/X vssd1 vssd1 vccd1 vccd1 _9787_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5066_ _9807_/Q vssd1 vssd1 vccd1 vccd1 _6317_/A sky130_fd_sc_hd__inv_2
XFILLER_84_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9874_ _9874_/CLK _9874_/D vssd1 vssd1 vccd1 vccd1 _9874_/Q sky130_fd_sc_hd__dfxtp_1
X_8825_ _8901_/C _8824_/A _8865_/C _8824_/Y vssd1 vssd1 vccd1 vccd1 _8825_/X sky130_fd_sc_hd__a22o_1
XFILLER_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8756_ _5858_/X _8754_/Y _8755_/X vssd1 vssd1 vccd1 vccd1 _8756_/Y sky130_fd_sc_hd__a21oi_1
X_5968_ _8008_/B vssd1 vssd1 vccd1 vccd1 _9503_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_12_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7707_ _7707_/A vssd1 vssd1 vccd1 vccd1 _7807_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4919_ _9868_/Q _4914_/X _9720_/Q _4912_/X _4915_/X vssd1 vssd1 vccd1 vccd1 _9868_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_178_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8687_ _8755_/A vssd1 vssd1 vccd1 vccd1 _8944_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_165_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5899_ _5903_/A _9141_/X vssd1 vssd1 vccd1 vccd1 _9610_/D sky130_fd_sc_hd__and2_1
XFILLER_165_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7638_ _7638_/A _7640_/B vssd1 vssd1 vccd1 vccd1 _7638_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7569_ _7470_/A _7470_/B _7470_/Y vssd1 vssd1 vccd1 vccd1 _7585_/A sky130_fd_sc_hd__o21ai_2
X_9308_ _9773_/Q _9307_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9308_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9239_ _7792_/Y _9752_/Q _9327_/S vssd1 vssd1 vccd1 vccd1 _9239_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6940_ _6903_/A _6903_/B _6925_/B vssd1 vssd1 vccd1 vccd1 _6941_/B sky130_fd_sc_hd__a21o_1
XFILLER_207_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6871_ _6872_/B _6881_/B vssd1 vssd1 vccd1 vccd1 _6877_/C sky130_fd_sc_hd__nor2_1
XFILLER_62_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8610_ _8823_/A _8610_/B _8610_/C vssd1 vssd1 vccd1 vccd1 _8611_/A sky130_fd_sc_hd__and3_1
X_9590_ _9836_/CLK _9590_/D vssd1 vssd1 vccd1 vccd1 _9590_/Q sky130_fd_sc_hd__dfxtp_1
X_5822_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5822_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_210_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8541_ _8498_/X _8513_/X _8481_/X _8514_/X vssd1 vssd1 vccd1 vccd1 _8541_/X sky130_fd_sc_hd__o22a_1
XFILLER_179_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5753_ _5721_/X _5722_/Y _5723_/X _5752_/X vssd1 vssd1 vccd1 vccd1 _5753_/X sky130_fd_sc_hd__o22a_1
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8472_ _8472_/A _9379_/X _8472_/C vssd1 vssd1 vccd1 vccd1 _8472_/X sky130_fd_sc_hd__or3_4
XFILLER_147_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5684_ _5692_/A vssd1 vssd1 vccd1 vccd1 _5684_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7423_ _7397_/X _7400_/X _7401_/X _7422_/X _7381_/X vssd1 vssd1 vccd1 vccd1 _7423_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_162_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7354_ _7327_/X _7331_/X _7332_/X _7353_/X _7311_/X vssd1 vssd1 vccd1 vccd1 _7354_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_190_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6305_ _9782_/Q vssd1 vssd1 vccd1 vccd1 _6487_/A sky130_fd_sc_hd__inv_2
XFILLER_116_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9024_ _9786_/Q _9903_/Q _9480_/S vssd1 vssd1 vccd1 vccd1 _9024_/X sky130_fd_sc_hd__mux2_1
X_7285_ _7311_/A _9471_/X _7331_/A _9472_/X vssd1 vssd1 vccd1 vccd1 _7286_/A sky130_fd_sc_hd__o22a_1
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6236_ _9582_/Q vssd1 vssd1 vccd1 vccd1 _8019_/A sky130_fd_sc_hd__inv_2
XFILLER_103_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6167_ _6167_/A vssd1 vssd1 vccd1 vccd1 _6168_/A sky130_fd_sc_hd__clkbuf_4
X_5118_ _9828_/Q vssd1 vssd1 vccd1 vccd1 _5118_/Y sky130_fd_sc_hd__inv_2
X_6098_ _7995_/A _9647_/Q _6088_/A _6085_/X vssd1 vssd1 vccd1 vccd1 _6098_/X sky130_fd_sc_hd__o22a_1
XFILLER_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9926_ _9926_/CLK _9926_/D vssd1 vssd1 vccd1 vccd1 _9926_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_150_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5049_ _5138_/A _9528_/Q vssd1 vssd1 vccd1 vccd1 _5097_/A sky130_fd_sc_hd__or2_4
XFILLER_198_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9857_ _9858_/CLK _9857_/D vssd1 vssd1 vccd1 vccd1 _9857_/Q sky130_fd_sc_hd__dfxtp_1
X_8808_ _8806_/Y _8807_/X _8806_/Y _8807_/X vssd1 vssd1 vccd1 vccd1 _8808_/X sky130_fd_sc_hd__o2bb2a_2
X_9788_ _9819_/CLK _9788_/D vssd1 vssd1 vccd1 vccd1 _9788_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_25_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8739_ _8732_/X _8738_/X _8732_/X _8738_/X vssd1 vssd1 vccd1 vccd1 _8739_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_139_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _9697_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _9887_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7070_ _7070_/A _7070_/B vssd1 vssd1 vccd1 vccd1 _7071_/B sky130_fd_sc_hd__or2_1
XFILLER_140_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6021_ _7947_/A _9639_/Q _6008_/A _6006_/X vssd1 vssd1 vccd1 vccd1 _6021_/X sky130_fd_sc_hd__o22a_1
XFILLER_82_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7972_ _8010_/B vssd1 vssd1 vccd1 vccd1 _7993_/B sky130_fd_sc_hd__clkbuf_2
X_9711_ _9828_/CLK _9711_/D vssd1 vssd1 vccd1 vccd1 _9711_/Q sky130_fd_sc_hd__dfxtp_1
X_6923_ _6859_/B _6922_/Y _6859_/B _6922_/Y vssd1 vssd1 vccd1 vccd1 _6923_/Y sky130_fd_sc_hd__a2bb2oi_2
XFILLER_207_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9642_ _9828_/CLK _9642_/D vssd1 vssd1 vccd1 vccd1 _9642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6854_ _6790_/X _6837_/X _6838_/X _6853_/X vssd1 vssd1 vccd1 vccd1 _6857_/A sky130_fd_sc_hd__o22a_1
XPHY_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5805_ _9654_/Q _5793_/X _5787_/X _7085_/A _5791_/X vssd1 vssd1 vccd1 vccd1 _9654_/D
+ sky130_fd_sc_hd__o221a_1
X_9573_ _9888_/CLK _9573_/D vssd1 vssd1 vccd1 vccd1 _9573_/Q sky130_fd_sc_hd__dfxtp_1
X_6785_ _6785_/A _6785_/B vssd1 vssd1 vccd1 vccd1 _6786_/B sky130_fd_sc_hd__or2_2
XFILLER_210_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8524_ _8390_/X _8402_/X _8390_/X _8402_/X vssd1 vssd1 vccd1 vccd1 _8525_/A sky130_fd_sc_hd__a2bb2o_1
X_5736_ _6556_/A _9656_/Q _5734_/A _5735_/Y vssd1 vssd1 vccd1 vccd1 _5736_/X sky130_fd_sc_hd__a22o_1
X_8455_ _8455_/A _8455_/B vssd1 vssd1 vccd1 vccd1 _8455_/Y sky130_fd_sc_hd__nor2_2
X_5667_ _9670_/Q vssd1 vssd1 vccd1 vccd1 _6569_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_129_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7406_ _7393_/X _7394_/X _7393_/X _7394_/X vssd1 vssd1 vccd1 vccd1 _7406_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_209_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5598_ _5609_/A _5598_/B vssd1 vssd1 vccd1 vccd1 _9706_/D sky130_fd_sc_hd__nor2_1
X_8386_ _9693_/Q _8386_/B vssd1 vssd1 vccd1 vccd1 _8386_/Y sky130_fd_sc_hd__nor2_1
XFILLER_190_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7337_ _7331_/C _7336_/A _7330_/A _7336_/Y vssd1 vssd1 vccd1 vccd1 _7337_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7268_ _7317_/A _9469_/X vssd1 vssd1 vccd1 vccd1 _7268_/X sky130_fd_sc_hd__or2_1
X_9007_ _9781_/Q _9898_/Q _9480_/S vssd1 vssd1 vccd1 vccd1 _9007_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6219_ _9579_/Q vssd1 vssd1 vccd1 vccd1 _8013_/A sky130_fd_sc_hd__inv_2
XINSDIODE2_10 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7199_ _7497_/A _7491_/B _7201_/A _9415_/X vssd1 vssd1 vccd1 vccd1 _7200_/B sky130_fd_sc_hd__o22a_1
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9909_ _9909_/CLK _9909_/D vssd1 vssd1 vccd1 vccd1 _9909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6570_ _6569_/A _6553_/B _6554_/B vssd1 vssd1 vccd1 vccd1 _6570_/X sky130_fd_sc_hd__a21bo_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5521_ _9490_/X _5510_/X _5621_/A vssd1 vssd1 vccd1 vccd1 _5617_/A sky130_fd_sc_hd__o21ai_1
XFILLER_145_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8240_ _9758_/Q _8240_/B vssd1 vssd1 vccd1 vccd1 _8240_/X sky130_fd_sc_hd__or2_1
XFILLER_172_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5452_ _9347_/X _9345_/X _5434_/Y _5507_/A vssd1 vssd1 vccd1 vccd1 _5503_/A sky130_fd_sc_hd__o22a_1
X_8171_ _7683_/A _8094_/X _7684_/A _8091_/X _8170_/X vssd1 vssd1 vccd1 vccd1 _8171_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_172_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5383_ _5383_/A vssd1 vssd1 vccd1 vccd1 _9722_/D sky130_fd_sc_hd__inv_2
XFILLER_125_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7122_ _7121_/A _7121_/B _7121_/X vssd1 vssd1 vccd1 vccd1 _7122_/X sky130_fd_sc_hd__a21bo_1
X_7053_ _6678_/A _6867_/B _6573_/X _6683_/A vssd1 vssd1 vccd1 vccd1 _7054_/B sky130_fd_sc_hd__o22a_1
XFILLER_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6004_ _9639_/Q vssd1 vssd1 vccd1 vccd1 _6004_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7955_ _7955_/A _7981_/B vssd1 vssd1 vccd1 vccd1 _7955_/X sky130_fd_sc_hd__or2_1
XFILLER_54_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7886_ _7885_/X _7879_/Y _7681_/B vssd1 vssd1 vccd1 vccd1 _7886_/Y sky130_fd_sc_hd__o21ai_1
X_6906_ _6880_/X _6883_/X _6884_/X _6905_/X _6864_/X vssd1 vssd1 vccd1 vccd1 _6906_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9625_ _9715_/CLK _9625_/D vssd1 vssd1 vccd1 vccd1 _9625_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_23_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6837_ _6810_/X _6814_/X _6815_/X _6836_/X _6794_/X vssd1 vssd1 vccd1 vccd1 _6837_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_210_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9556_ _9924_/CLK _9556_/D vssd1 vssd1 vccd1 vccd1 _9556_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8507_ _8505_/X _8506_/Y _8505_/X _8506_/Y vssd1 vssd1 vccd1 vccd1 _8508_/A sky130_fd_sc_hd__a2bb2o_1
X_6768_ _6812_/A _9094_/X _6814_/A _9095_/X vssd1 vssd1 vccd1 vccd1 _6769_/A sky130_fd_sc_hd__o22a_1
XFILLER_50_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5719_ _9679_/Q _9662_/Q _5717_/Y _5718_/Y vssd1 vssd1 vccd1 vccd1 _5719_/X sky130_fd_sc_hd__a22o_1
X_9487_ _9486_/X _8959_/A _9505_/S vssd1 vssd1 vccd1 vccd1 _9487_/X sky130_fd_sc_hd__mux2_1
X_6699_ _6971_/A _6766_/B _7005_/A _6721_/B vssd1 vssd1 vccd1 vccd1 _6701_/A sky130_fd_sc_hd__o22a_1
XFILLER_40_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8438_ _8472_/C _8438_/B vssd1 vssd1 vccd1 vccd1 _8460_/A sky130_fd_sc_hd__nand2_4
XFILLER_163_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8369_ _8369_/A _8369_/B _8369_/C _8369_/D vssd1 vssd1 vccd1 vccd1 _8374_/A sky130_fd_sc_hd__and4_1
XFILLER_136_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput6 io_wb_adr_i[1] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7740_ _7895_/A _8200_/A _4843_/X _6360_/Y _7739_/X vssd1 vssd1 vccd1 vccd1 _7752_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_91_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4952_ _4952_/A vssd1 vssd1 vccd1 vccd1 _4952_/X sky130_fd_sc_hd__buf_1
X_7671_ _9914_/Q _7671_/B vssd1 vssd1 vccd1 vccd1 _7846_/A sky130_fd_sc_hd__or2_1
X_4883_ _9739_/Q _4879_/X _9887_/Q _4880_/X _4881_/X vssd1 vssd1 vccd1 vccd1 _9887_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_189_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6622_ _6622_/A _6622_/B vssd1 vssd1 vccd1 vccd1 _6622_/Y sky130_fd_sc_hd__nor2_1
X_9410_ _8008_/X _6110_/Y _9504_/S vssd1 vssd1 vccd1 vccd1 _9410_/X sky130_fd_sc_hd__mux2_1
X_6553_ _6569_/A _6553_/B vssd1 vssd1 vccd1 vccd1 _6554_/B sky130_fd_sc_hd__or2_1
X_9341_ _7051_/Y _7628_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9341_/X sky130_fd_sc_hd__mux2_1
X_6484_ _6487_/A _6487_/B _6304_/Y _6482_/X vssd1 vssd1 vccd1 vccd1 _6494_/A sky130_fd_sc_hd__o22a_1
XFILLER_145_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9272_ _9760_/Q _9271_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9272_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5504_ _5431_/A _5431_/B _5431_/Y vssd1 vssd1 vccd1 vccd1 _5504_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_145_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8223_ _8223_/A _8227_/B vssd1 vssd1 vccd1 vccd1 _8223_/Y sky130_fd_sc_hd__nor2_1
X_5435_ _9354_/X _9352_/X _9354_/X _9352_/X vssd1 vssd1 vccd1 vccd1 _5435_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8154_ _7743_/A _8109_/X _8153_/Y vssd1 vssd1 vccd1 vccd1 _8154_/Y sky130_fd_sc_hd__o21bai_1
X_5366_ _5366_/A vssd1 vssd1 vccd1 vccd1 _9726_/D sky130_fd_sc_hd__inv_2
X_8085_ _9557_/Q _8085_/B vssd1 vssd1 vccd1 vccd1 _8093_/A sky130_fd_sc_hd__or2_1
XFILLER_141_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5297_ _5297_/A vssd1 vssd1 vccd1 vccd1 _9737_/D sky130_fd_sc_hd__inv_2
X_7105_ _7156_/A vssd1 vssd1 vccd1 vccd1 _7487_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_59_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7036_ _7010_/X _7011_/X _7012_/X _7035_/X vssd1 vssd1 vccd1 vccd1 _7036_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_101_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8987_ _7990_/X _6074_/B _9504_/S vssd1 vssd1 vccd1 vccd1 _8987_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7938_ _8472_/A vssd1 vssd1 vccd1 vccd1 _8576_/A sky130_fd_sc_hd__buf_1
XFILLER_82_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7869_ _7869_/A _7869_/B vssd1 vssd1 vccd1 vccd1 _7873_/B sky130_fd_sc_hd__or2_2
XPHY_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9608_ _9895_/CLK _9608_/D vssd1 vssd1 vccd1 vccd1 _9608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9539_ _9907_/CLK _9539_/D vssd1 vssd1 vccd1 vccd1 _9539_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5220_ _5041_/X _5151_/X _9748_/Q _5152_/X _5214_/X vssd1 vssd1 vccd1 vccd1 _9748_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5151_ _5203_/A vssd1 vssd1 vccd1 vccd1 _5151_/X sky130_fd_sc_hd__buf_2
XFILLER_130_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5082_ _5061_/X _6317_/D _5081_/Y _5073_/X vssd1 vssd1 vccd1 vccd1 _5083_/B sky130_fd_sc_hd__o22a_1
XFILLER_96_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8910_ _8938_/A _8942_/B _8944_/C _9419_/X vssd1 vssd1 vccd1 vccd1 _8910_/X sky130_fd_sc_hd__o22a_1
XFILLER_96_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9890_ _9893_/CLK _9890_/D vssd1 vssd1 vccd1 vccd1 _9890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8841_ _8841_/A _8841_/B vssd1 vssd1 vccd1 vccd1 _8887_/A sky130_fd_sc_hd__or2_1
X_8772_ _8800_/A _8773_/D _8773_/C _8725_/B vssd1 vssd1 vccd1 vccd1 _8775_/A sky130_fd_sc_hd__o22a_1
XFILLER_92_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7723_ _7723_/A vssd1 vssd1 vccd1 vccd1 _7723_/X sky130_fd_sc_hd__clkbuf_2
X_5984_ _9850_/Q vssd1 vssd1 vccd1 vccd1 _7935_/A sky130_fd_sc_hd__inv_2
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4935_ _4952_/A vssd1 vssd1 vccd1 vccd1 _4935_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_177_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7654_ _9901_/Q vssd1 vssd1 vccd1 vccd1 _7793_/A sky130_fd_sc_hd__inv_2
X_4866_ _4880_/A vssd1 vssd1 vccd1 vccd1 _4866_/X sky130_fd_sc_hd__buf_1
XFILLER_177_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4797_ _9918_/Q vssd1 vssd1 vccd1 vccd1 _4798_/A sky130_fd_sc_hd__clkbuf_2
X_6605_ _6872_/B vssd1 vssd1 vccd1 vccd1 _6868_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7585_ _7585_/A vssd1 vssd1 vccd1 vccd1 _7597_/A sky130_fd_sc_hd__inv_2
X_9324_ _9777_/Q _9323_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9324_/X sky130_fd_sc_hd__mux2_1
X_6536_ _6542_/A vssd1 vssd1 vccd1 vccd1 _6541_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6467_ _6467_/A vssd1 vssd1 vccd1 vccd1 _6467_/Y sky130_fd_sc_hd__inv_2
X_9255_ _7809_/Y _9756_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9255_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6398_ _6354_/Y _6397_/Y _9779_/Q _6397_/A vssd1 vssd1 vccd1 vccd1 _6550_/B sky130_fd_sc_hd__o22a_1
X_8206_ _5162_/X _8205_/X _8200_/B vssd1 vssd1 vccd1 vccd1 _8206_/X sky130_fd_sc_hd__a21bo_1
XFILLER_133_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9186_ _6527_/Y _9791_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9540_/D sky130_fd_sc_hd__mux2_1
X_5418_ _5418_/A _5418_/B vssd1 vssd1 vccd1 vccd1 _5418_/Y sky130_fd_sc_hd__nor2_1
X_8137_ _9901_/Q _8124_/X _9902_/Q _8123_/B _8136_/X vssd1 vssd1 vccd1 vccd1 _8137_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_121_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5349_ _5363_/A vssd1 vssd1 vccd1 vccd1 _5349_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8068_ _9540_/Q _8068_/B vssd1 vssd1 vccd1 vccd1 _8069_/B sky130_fd_sc_hd__or2_1
X_7019_ _6920_/X _6959_/X _6920_/X _6959_/X vssd1 vssd1 vccd1 vccd1 _7019_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput31 io_wb_dat_i[23] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_4
Xinput20 io_wb_dat_i[13] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_4
XFILLER_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput42 io_wb_dat_i[4] vssd1 vssd1 vccd1 vccd1 _4978_/A sky130_fd_sc_hd__buf_6
X_7370_ _7356_/X _7357_/X _7358_/X _7369_/X vssd1 vssd1 vccd1 vccd1 _7370_/X sky130_fd_sc_hd__o22a_1
X_6321_ _6542_/A vssd1 vssd1 vccd1 vccd1 _9178_/S sky130_fd_sc_hd__inv_2
XFILLER_155_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6252_ _9583_/Q _6171_/X _6243_/A _6248_/A vssd1 vssd1 vccd1 vccd1 _6252_/X sky130_fd_sc_hd__a22o_1
XFILLER_143_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9040_ _7992_/Y _9039_/X _9052_/S vssd1 vssd1 vccd1 vccd1 _9040_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5203_ _5203_/A vssd1 vssd1 vccd1 vccd1 _5203_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6183_ _7976_/A _6143_/X _6187_/A vssd1 vssd1 vccd1 vccd1 _6183_/Y sky130_fd_sc_hd__o21ai_1
X_5134_ _5128_/X _9788_/Q _5130_/X _9215_/X _5132_/X vssd1 vssd1 vccd1 vccd1 _9788_/D
+ sky130_fd_sc_hd__o221a_1
X_5065_ _5069_/A _5065_/B vssd1 vssd1 vccd1 vccd1 _9808_/D sky130_fd_sc_hd__nor2_1
XFILLER_111_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9873_ _9874_/CLK _9873_/D vssd1 vssd1 vccd1 vccd1 _9873_/Q sky130_fd_sc_hd__dfxtp_1
X_8824_ _8824_/A vssd1 vssd1 vccd1 vccd1 _8824_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8755_ _8755_/A _9396_/X vssd1 vssd1 vccd1 vccd1 _8755_/X sky130_fd_sc_hd__or2_1
X_5967_ _5967_/A vssd1 vssd1 vccd1 vccd1 _8008_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_178_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8686_ _8686_/A vssd1 vssd1 vccd1 vccd1 _8735_/C sky130_fd_sc_hd__inv_2
X_7706_ _9904_/Q vssd1 vssd1 vccd1 vccd1 _7707_/A sky130_fd_sc_hd__inv_2
X_4918_ _9869_/Q _4914_/X _9721_/Q _4912_/X _4915_/X vssd1 vssd1 vccd1 vccd1 _9869_/D
+ sky130_fd_sc_hd__o221a_1
X_7637_ _7637_/A _7640_/B vssd1 vssd1 vccd1 vccd1 _7637_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5898_ _5910_/A vssd1 vssd1 vccd1 vccd1 _5903_/A sky130_fd_sc_hd__buf_1
X_4849_ _9898_/Q vssd1 vssd1 vccd1 vccd1 _7749_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_148_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7568_ _7548_/A _7548_/B _7548_/X vssd1 vssd1 vccd1 vccd1 _7584_/A sky130_fd_sc_hd__a21bo_1
XFILLER_180_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9307_ _7880_/X _9773_/Q _9327_/S vssd1 vssd1 vccd1 vccd1 _9307_/X sky130_fd_sc_hd__mux2_1
X_6519_ _6522_/A _6519_/B vssd1 vssd1 vccd1 vccd1 _6519_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7499_ _7487_/A _9432_/X _7518_/A _7491_/B vssd1 vssd1 vccd1 vccd1 _7500_/B sky130_fd_sc_hd__o22a_1
XFILLER_161_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9238_ _9237_/X _5035_/A _9306_/S vssd1 vssd1 vccd1 vccd1 _9238_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9169_ _6298_/Y input39/X _9170_/S vssd1 vssd1 vccd1 vccd1 _9169_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6870_ _6868_/X _6869_/X _6868_/X _6869_/X vssd1 vssd1 vccd1 vccd1 _6876_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5821_ _9649_/Q _5818_/X input21/X _5819_/X _5809_/X vssd1 vssd1 vccd1 vccd1 _9649_/D
+ sky130_fd_sc_hd__o221a_1
X_8540_ _8533_/X _8539_/X _8533_/X _8539_/X vssd1 vssd1 vccd1 vccd1 _8540_/X sky130_fd_sc_hd__a2bb2o_1
X_5752_ _8386_/B _5726_/Y _5727_/X _5751_/X vssd1 vssd1 vccd1 vccd1 _5752_/X sky130_fd_sc_hd__o22a_1
XFILLER_203_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8471_ _8471_/A _9377_/X vssd1 vssd1 vccd1 vccd1 _8576_/C sky130_fd_sc_hd__or2_4
X_5683_ _6578_/A _5681_/X _9106_/X _5676_/X _5682_/X vssd1 vssd1 vccd1 vccd1 _9679_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7422_ _7416_/A _7443_/A _7415_/Y _7413_/A _7421_/Y vssd1 vssd1 vccd1 vccd1 _7422_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_162_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7353_ _7351_/A _7348_/X _7350_/X _7352_/Y vssd1 vssd1 vccd1 vccd1 _7353_/X sky130_fd_sc_hd__o22a_1
XFILLER_190_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6304_ _9783_/Q vssd1 vssd1 vccd1 vccd1 _6304_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_2_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _9917_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_103_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7284_ _7280_/X _7283_/X _7280_/X _7283_/X vssd1 vssd1 vccd1 vccd1 _7284_/X sky130_fd_sc_hd__a2bb2o_1
X_9023_ _7957_/Y _9600_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9023_/X sky130_fd_sc_hd__mux2_1
X_6235_ _6244_/A _6234_/X _6244_/A _6234_/X vssd1 vssd1 vccd1 vccd1 _6235_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6166_ _6166_/A vssd1 vssd1 vccd1 vccd1 _6167_/A sky130_fd_sc_hd__clkbuf_2
X_5117_ _9796_/Q vssd1 vssd1 vccd1 vccd1 _6500_/A sky130_fd_sc_hd__inv_2
X_6097_ _6095_/X _6096_/Y _6095_/X _6096_/Y vssd1 vssd1 vccd1 vccd1 _6097_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9925_ _9926_/CLK _9925_/D vssd1 vssd1 vccd1 vccd1 _9925_/Q sky130_fd_sc_hd__dfxtp_1
X_5048_ _5048_/A vssd1 vssd1 vccd1 vccd1 _5138_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9856_ _9858_/CLK _9856_/D vssd1 vssd1 vccd1 vccd1 _9856_/Q sky130_fd_sc_hd__dfxtp_2
X_8807_ _8807_/A _8893_/B _8807_/C vssd1 vssd1 vccd1 vccd1 _8807_/X sky130_fd_sc_hd__or3_1
X_9787_ _9929_/CLK _9787_/D vssd1 vssd1 vccd1 vccd1 _9787_/Q sky130_fd_sc_hd__dfxtp_1
X_8738_ _8823_/C _8737_/B _8762_/A vssd1 vssd1 vccd1 vccd1 _8738_/X sky130_fd_sc_hd__a21bo_1
X_6999_ _6995_/X _6996_/X _6995_/X _6996_/X vssd1 vssd1 vccd1 vccd1 _7003_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8669_ _8766_/C vssd1 vssd1 vccd1 vccd1 _8712_/C sky130_fd_sc_hd__inv_2
XFILLER_178_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6020_ _6019_/A _6018_/Y _6019_/Y _6018_/A vssd1 vssd1 vccd1 vccd1 _6020_/X sky130_fd_sc_hd__o22a_1
XFILLER_67_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7971_ _7971_/A vssd1 vssd1 vccd1 vccd1 _8010_/B sky130_fd_sc_hd__buf_1
X_9710_ _9828_/CLK _9710_/D vssd1 vssd1 vccd1 vccd1 _9710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6922_ _6777_/X _6855_/Y _6859_/A vssd1 vssd1 vccd1 vccd1 _6922_/Y sky130_fd_sc_hd__o21ai_2
X_9641_ _9828_/CLK _9641_/D vssd1 vssd1 vccd1 vccd1 _9641_/Q sky130_fd_sc_hd__dfxtp_1
X_6853_ _6839_/X _6840_/X _6841_/X _6852_/X vssd1 vssd1 vccd1 vccd1 _6853_/X sky130_fd_sc_hd__o22a_1
X_5804_ _5745_/X _5803_/X _5745_/X _5803_/X vssd1 vssd1 vccd1 vccd1 _7085_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_200_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6784_ _6760_/C _6757_/B _6757_/Y vssd1 vssd1 vccd1 vccd1 _6785_/B sky130_fd_sc_hd__o21ai_2
XFILLER_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9572_ _9578_/CLK _9572_/D vssd1 vssd1 vccd1 vccd1 _9572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8523_ _8522_/A _8522_/B _8555_/A vssd1 vssd1 vccd1 vccd1 _8523_/X sky130_fd_sc_hd__a21bo_1
X_5735_ _9656_/Q vssd1 vssd1 vccd1 vccd1 _5735_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8454_ _8452_/X _8453_/Y _8452_/X _8453_/Y vssd1 vssd1 vccd1 vccd1 _8455_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5666_ _9687_/Q _5658_/X _8394_/B _5662_/X _5660_/X vssd1 vssd1 vccd1 vccd1 _9687_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_108_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7405_ _7405_/A _7405_/B vssd1 vssd1 vccd1 vccd1 _7416_/A sky130_fd_sc_hd__or2_1
X_5597_ _5586_/X _5594_/Y _5595_/Y _7643_/A _5577_/X vssd1 vssd1 vccd1 vccd1 _5598_/B
+ sky130_fd_sc_hd__o32a_1
X_8385_ _9694_/Q _5721_/X _9694_/Q _5721_/X vssd1 vssd1 vccd1 vccd1 _8385_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_209_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7336_ _7336_/A vssd1 vssd1 vccd1 vccd1 _7336_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7267_ _7311_/A _9471_/X _7331_/A _9472_/X vssd1 vssd1 vccd1 vccd1 _7267_/X sky130_fd_sc_hd__or4_4
X_9006_ _9005_/X _9595_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9006_/X sky130_fd_sc_hd__mux2_1
X_6218_ _6221_/D _6217_/Y _6221_/D _6217_/Y vssd1 vssd1 vccd1 vccd1 _6218_/X sky130_fd_sc_hd__a2bb2o_1
X_7198_ _9414_/X vssd1 vssd1 vccd1 vccd1 _7491_/B sky130_fd_sc_hd__buf_1
XFILLER_58_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_11 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6149_ _9567_/Q _6165_/A _7949_/A _6148_/X vssd1 vssd1 vccd1 vccd1 _6152_/A sky130_fd_sc_hd__a22o_1
X_9908_ _9909_/CLK _9908_/D vssd1 vssd1 vccd1 vccd1 _9908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9839_ _9898_/CLK _9839_/D vssd1 vssd1 vccd1 vccd1 _9839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5520_ _5626_/A _5622_/B vssd1 vssd1 vccd1 vccd1 _5621_/A sky130_fd_sc_hd__or2_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5451_ _9354_/X _9352_/X _5435_/X _5450_/X vssd1 vssd1 vccd1 vccd1 _5507_/A sky130_fd_sc_hd__o22a_1
X_8170_ _4775_/X _8095_/Y _7683_/A _8094_/X _8169_/X vssd1 vssd1 vccd1 vccd1 _8170_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5382_ _5376_/B _5379_/X _5381_/Y _5329_/A _5364_/X vssd1 vssd1 vccd1 vccd1 _5383_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_172_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7121_ _7121_/A _7121_/B vssd1 vssd1 vccd1 vccd1 _7121_/X sky130_fd_sc_hd__or2_1
XFILLER_99_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7052_ _6833_/A _6833_/B _6834_/B vssd1 vssd1 vccd1 vccd1 _7069_/A sky130_fd_sc_hd__a21bo_1
X_6003_ _9852_/Q vssd1 vssd1 vccd1 vccd1 _7947_/A sky130_fd_sc_hd__inv_2
XFILLER_86_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7954_ _8008_/B vssd1 vssd1 vccd1 vccd1 _7981_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6905_ _6899_/A _6926_/A _6898_/Y _6896_/A _6904_/Y vssd1 vssd1 vccd1 vccd1 _6905_/X
+ sky130_fd_sc_hd__o32a_1
XPHY_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7885_ _7887_/A vssd1 vssd1 vccd1 vccd1 _7885_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_20_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _9699_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6836_ _6830_/A _6847_/A _6829_/Y _6827_/A _6835_/Y vssd1 vssd1 vccd1 vccd1 _6836_/X
+ sky130_fd_sc_hd__o32a_1
X_9624_ _9858_/CLK _9624_/D vssd1 vssd1 vccd1 vccd1 _9624_/Q sky130_fd_sc_hd__dfxtp_1
X_9555_ _9924_/CLK _9555_/D vssd1 vssd1 vccd1 vccd1 _9555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6767_ _6763_/X _6766_/X _6763_/X _6766_/X vssd1 vssd1 vccd1 vccd1 _6767_/X sky130_fd_sc_hd__a2bb2o_1
X_8506_ _8475_/C _8455_/Y _9628_/Q _8500_/Y vssd1 vssd1 vccd1 vccd1 _8506_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_183_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5718_ _9662_/Q vssd1 vssd1 vccd1 vccd1 _5718_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9486_ _7947_/X _6004_/Y _9504_/S vssd1 vssd1 vccd1 vccd1 _9486_/X sky130_fd_sc_hd__mux2_1
X_6698_ _6764_/B vssd1 vssd1 vccd1 vccd1 _6721_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_35_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _9893_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8437_ _8475_/C _8436_/X _8475_/C _8436_/X vssd1 vssd1 vccd1 vccd1 _8438_/B sky130_fd_sc_hd__o2bb2a_2
XFILLER_163_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5649_ _9677_/Q vssd1 vssd1 vccd1 vccd1 _6576_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8368_ _4765_/A _8088_/Y _8357_/A _8367_/X vssd1 vssd1 vccd1 vccd1 _8368_/X sky130_fd_sc_hd__o22a_1
XFILLER_156_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7319_ _7321_/B vssd1 vssd1 vccd1 vccd1 _7408_/B sky130_fd_sc_hd__clkbuf_2
X_8299_ _6354_/Y _8209_/Y _6550_/B _8199_/B vssd1 vssd1 vccd1 vccd1 _8301_/B sky130_fd_sc_hd__o22a_1
XFILLER_104_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 io_wb_adr_i[2] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4951_ _4951_/A vssd1 vssd1 vccd1 vccd1 _4951_/X sky130_fd_sc_hd__buf_1
X_7670_ _9913_/Q _7837_/A vssd1 vssd1 vccd1 vccd1 _7671_/B sky130_fd_sc_hd__or2_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4882_ _9740_/Q _4879_/X _9888_/Q _4880_/X _4881_/X vssd1 vssd1 vccd1 vccd1 _9888_/D
+ sky130_fd_sc_hd__a221o_1
X_6621_ _7006_/A _6971_/B _6691_/C vssd1 vssd1 vccd1 vccd1 _6622_/B sky130_fd_sc_hd__or3_1
XFILLER_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9340_ _7607_/X _7578_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9340_/X sky130_fd_sc_hd__mux2_4
XFILLER_158_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6552_ _6571_/A _6804_/C vssd1 vssd1 vccd1 vccd1 _6553_/B sky130_fd_sc_hd__or2_1
XFILLER_173_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6483_ _8056_/A _5218_/X _6367_/A _6327_/Y _6367_/Y vssd1 vssd1 vccd1 vccd1 _6487_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_118_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9271_ _7826_/Y _9760_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9271_/X sky130_fd_sc_hd__mux2_1
X_5503_ _5503_/A vssd1 vssd1 vccd1 vccd1 _5503_/Y sky130_fd_sc_hd__inv_2
X_8222_ _6351_/A _8221_/X _8219_/X vssd1 vssd1 vccd1 vccd1 _8222_/X sky130_fd_sc_hd__a21bo_1
XFILLER_106_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5434_ _5434_/A _5434_/B vssd1 vssd1 vccd1 vccd1 _5434_/Y sky130_fd_sc_hd__nor2_1
XFILLER_145_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8153_ _7743_/A _8109_/X _7715_/X _8110_/X _8152_/X vssd1 vssd1 vccd1 vccd1 _8153_/Y
+ sky130_fd_sc_hd__a221oi_2
XFILLER_10_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5365_ _5358_/B _5356_/X _5362_/Y _5333_/A _5364_/X vssd1 vssd1 vccd1 vccd1 _5366_/A
+ sky130_fd_sc_hd__o32a_1
X_7104_ _7324_/A vssd1 vssd1 vccd1 vccd1 _7156_/A sky130_fd_sc_hd__clkbuf_2
X_8084_ _9556_/Q _8084_/B vssd1 vssd1 vccd1 vccd1 _8085_/B sky130_fd_sc_hd__or2_1
XFILLER_113_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5296_ _5291_/B _5224_/A _5295_/Y _5275_/A _5242_/A vssd1 vssd1 vccd1 vccd1 _5297_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7035_ _7013_/X _7014_/X _7015_/X _7034_/X vssd1 vssd1 vccd1 vccd1 _7035_/X sky130_fd_sc_hd__o22a_1
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8986_ _8985_/X _6337_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _8986_/X sky130_fd_sc_hd__mux2_2
XFILLER_82_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7937_ _9630_/Q vssd1 vssd1 vccd1 vccd1 _8472_/A sky130_fd_sc_hd__inv_2
XFILLER_42_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7868_ _7869_/A _7863_/Y _7677_/B vssd1 vssd1 vccd1 vccd1 _7868_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_23_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9607_ _9895_/CLK _9607_/D vssd1 vssd1 vccd1 vccd1 _9607_/Q sky130_fd_sc_hd__dfxtp_1
X_6819_ _6819_/A _6819_/B vssd1 vssd1 vccd1 vccd1 _6830_/A sky130_fd_sc_hd__or2_1
X_7799_ _7797_/A _7797_/B _7798_/Y _7790_/X vssd1 vssd1 vccd1 vccd1 _7799_/Y sky130_fd_sc_hd__a211oi_2
XPHY_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9538_ _9907_/CLK _9538_/D vssd1 vssd1 vccd1 vccd1 _9538_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9469_ _7090_/X _6118_/Y _9475_/S vssd1 vssd1 vccd1 vccd1 _9469_/X sky130_fd_sc_hd__mux2_4
XFILLER_136_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5150_ _5178_/A vssd1 vssd1 vccd1 vccd1 _5203_/A sky130_fd_sc_hd__buf_2
XFILLER_111_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5081_ _9836_/Q vssd1 vssd1 vccd1 vccd1 _5081_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8840_ _8840_/A vssd1 vssd1 vccd1 vccd1 _8841_/B sky130_fd_sc_hd__inv_2
XFILLER_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8771_ _8767_/X _8770_/X _8767_/X _8770_/X vssd1 vssd1 vccd1 vccd1 _8771_/X sky130_fd_sc_hd__a2bb2o_1
X_5983_ _9848_/Q _5703_/B _5981_/A _5704_/C _5981_/Y vssd1 vssd1 vccd1 vccd1 _5983_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_52_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7722_ _7848_/A vssd1 vssd1 vccd1 vccd1 _7723_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4934_ _4951_/A vssd1 vssd1 vccd1 vccd1 _4934_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_177_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7653_ _7776_/A vssd1 vssd1 vccd1 vccd1 _7778_/B sky130_fd_sc_hd__inv_2
X_4865_ _4879_/A vssd1 vssd1 vccd1 vccd1 _4865_/X sky130_fd_sc_hd__buf_1
XFILLER_60_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4796_ _4796_/A vssd1 vssd1 vccd1 vccd1 _4796_/X sky130_fd_sc_hd__buf_2
X_6604_ _9615_/Q vssd1 vssd1 vccd1 vccd1 _6872_/B sky130_fd_sc_hd__inv_2
X_7584_ _7584_/A vssd1 vssd1 vccd1 vccd1 _7598_/A sky130_fd_sc_hd__inv_2
X_9323_ _7900_/X _9777_/Q _9327_/S vssd1 vssd1 vccd1 vccd1 _9323_/X sky130_fd_sc_hd__mux2_1
X_6535_ _6535_/A _6535_/B vssd1 vssd1 vccd1 vccd1 _6535_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9254_ _9253_/X _5026_/A _9306_/S vssd1 vssd1 vccd1 vccd1 _9254_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8205_ _8205_/A _8205_/B vssd1 vssd1 vccd1 vccd1 _8205_/X sky130_fd_sc_hd__or2_1
X_6466_ _6463_/X _6466_/B _6466_/C _6466_/D vssd1 vssd1 vccd1 vccd1 _6466_/Y sky130_fd_sc_hd__nand4b_4
X_6397_ _6397_/A vssd1 vssd1 vccd1 vccd1 _6397_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9185_ _6526_/Y _9790_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9539_/D sky130_fd_sc_hd__mux2_1
X_5417_ _9361_/X vssd1 vssd1 vccd1 vccd1 _5418_/B sky130_fd_sc_hd__inv_2
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8136_ _7657_/A _8126_/Y _9901_/Q _8124_/X _8135_/X vssd1 vssd1 vccd1 vccd1 _8136_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_121_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5348_ _5919_/A _5348_/B vssd1 vssd1 vccd1 vccd1 _5363_/A sky130_fd_sc_hd__or2_1
X_8067_ _9539_/Q _8067_/B vssd1 vssd1 vccd1 vccd1 _8068_/B sky130_fd_sc_hd__or2_1
X_7018_ _7016_/X _7017_/X _7016_/X _7017_/X vssd1 vssd1 vccd1 vccd1 _7018_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5279_ _9741_/Q _5279_/B vssd1 vssd1 vccd1 vccd1 _5279_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8969_ vssd1 vssd1 vccd1 vccd1 _8969_/HI _9222_/A1 sky130_fd_sc_hd__conb_1
XPHY_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput21 io_wb_dat_i[14] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_6
Xinput10 io_wb_adr_i[5] vssd1 vssd1 vccd1 vccd1 _5707_/A sky130_fd_sc_hd__buf_1
Xinput32 io_wb_dat_i[24] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_4
XFILLER_162_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6320_ _6308_/X _6310_/X _6315_/Y _6319_/X vssd1 vssd1 vccd1 vccd1 _6542_/A sky130_fd_sc_hd__o211a_2
Xinput43 io_wb_dat_i[5] vssd1 vssd1 vccd1 vccd1 _5032_/A sky130_fd_sc_hd__buf_6
X_6251_ _9584_/Q _6169_/A _8024_/A _6245_/A vssd1 vssd1 vccd1 vccd1 _6265_/B sky130_fd_sc_hd__a22o_1
XFILLER_143_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5202_ input47/X _5192_/X _9757_/Q _5193_/X _5194_/X vssd1 vssd1 vccd1 vccd1 _9757_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6182_ _9572_/Q _6166_/A _7983_/A _6197_/A vssd1 vssd1 vccd1 vccd1 _6187_/B sky130_fd_sc_hd__a22o_1
X_5133_ _5128_/X _9789_/Q _5130_/X _9216_/X _5132_/X vssd1 vssd1 vccd1 vccd1 _9789_/D
+ sky130_fd_sc_hd__o221a_1
X_5064_ _5061_/X _6316_/D _5063_/Y _5050_/X vssd1 vssd1 vccd1 vccd1 _5065_/B sky130_fd_sc_hd__o22a_1
X_9872_ _9893_/CLK _9872_/D vssd1 vssd1 vccd1 vccd1 _9872_/Q sky130_fd_sc_hd__dfxtp_1
X_8823_ _8823_/A _8823_/B _8823_/C vssd1 vssd1 vccd1 vccd1 _8824_/A sky130_fd_sc_hd__and3_1
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8754_ _8821_/B vssd1 vssd1 vccd1 vccd1 _8754_/Y sky130_fd_sc_hd__inv_2
X_5966_ _9073_/X _5937_/A _9563_/Q _5938_/A vssd1 vssd1 vccd1 vccd1 _9563_/D sky130_fd_sc_hd__a22o_1
XFILLER_197_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8685_ _8751_/B vssd1 vssd1 vccd1 vccd1 _8823_/B sky130_fd_sc_hd__inv_2
X_7705_ _7705_/A _7705_/B _7705_/C _7705_/D vssd1 vssd1 vccd1 vccd1 _7773_/A sky130_fd_sc_hd__and4_1
X_5897_ _5041_/X _5884_/X _9611_/Q _5885_/X _5070_/A vssd1 vssd1 vccd1 vccd1 _9611_/D
+ sky130_fd_sc_hd__a221o_1
X_4917_ _9870_/Q _4914_/X _9722_/Q _4912_/X _4915_/X vssd1 vssd1 vccd1 vccd1 _9870_/D
+ sky130_fd_sc_hd__o221a_1
X_4848_ _9234_/X _4834_/X _4847_/X _4836_/X _4845_/X vssd1 vssd1 vccd1 vccd1 _9899_/D
+ sky130_fd_sc_hd__o221a_1
X_7636_ _7636_/A _7640_/B vssd1 vssd1 vccd1 vccd1 _7636_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4779_ _9322_/X _4763_/X _4775_/X _4767_/X _4778_/X vssd1 vssd1 vccd1 vccd1 _9925_/D
+ sky130_fd_sc_hd__o221a_1
X_9306_ _9305_/X input32/X _9306_/S vssd1 vssd1 vccd1 vccd1 _9306_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7567_ _7546_/X _7548_/X _7546_/X _7548_/X vssd1 vssd1 vccd1 vccd1 _7583_/A sky130_fd_sc_hd__a2bb2o_1
X_6518_ _6316_/A _6399_/Y _9178_/S _6517_/X vssd1 vssd1 vccd1 vccd1 _9206_/S sky130_fd_sc_hd__o211a_4
X_7498_ _7206_/X _7207_/X _7206_/X _7207_/X vssd1 vssd1 vccd1 vccd1 _7498_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_180_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9237_ _9236_/X _7791_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9237_/X sky130_fd_sc_hd__mux2_1
X_6449_ _6337_/A _6376_/B _6377_/B vssd1 vssd1 vccd1 vccd1 _6453_/B sky130_fd_sc_hd__a21bo_1
XFILLER_106_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9168_ _6293_/X input37/X _9170_/S vssd1 vssd1 vccd1 vccd1 _9168_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8119_ _9537_/Q _8065_/B _8066_/B vssd1 vssd1 vccd1 vccd1 _8119_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9099_ _6010_/Y _6011_/Y _9896_/Q vssd1 vssd1 vccd1 vccd1 _9099_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5820_ _9650_/Q _5818_/X input22/X _5819_/X _5809_/X vssd1 vssd1 vccd1 vccd1 _9650_/D
+ sky130_fd_sc_hd__o221a_1
X_5751_ _6582_/A _5729_/Y _5730_/X _5750_/X vssd1 vssd1 vccd1 vccd1 _5751_/X sky130_fd_sc_hd__o22a_1
XFILLER_34_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8470_ _8605_/A _9381_/X vssd1 vssd1 vccd1 vccd1 _8495_/A sky130_fd_sc_hd__or2_2
XFILLER_147_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5682_ _5772_/A vssd1 vssd1 vccd1 vccd1 _5682_/X sky130_fd_sc_hd__buf_1
X_7421_ _7421_/A _7442_/B vssd1 vssd1 vccd1 vccd1 _7421_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7352_ _7352_/A _7352_/B vssd1 vssd1 vccd1 vccd1 _7352_/Y sky130_fd_sc_hd__nor2_1
X_6303_ _8047_/B vssd1 vssd1 vccd1 vccd1 _8030_/B sky130_fd_sc_hd__clkbuf_4
X_7283_ _7491_/A _7283_/B _7283_/C vssd1 vssd1 vccd1 vccd1 _7283_/X sky130_fd_sc_hd__or3_1
X_9022_ _9021_/X _9753_/Q _9481_/S vssd1 vssd1 vccd1 vccd1 _9022_/X sky130_fd_sc_hd__mux2_2
X_6234_ _6244_/C _6234_/B vssd1 vssd1 vccd1 vccd1 _6234_/X sky130_fd_sc_hd__and2_1
XFILLER_116_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6165_ _6165_/A vssd1 vssd1 vccd1 vccd1 _6166_/A sky130_fd_sc_hd__clkbuf_2
X_5116_ _8177_/A vssd1 vssd1 vccd1 vccd1 _5579_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6096_ _9860_/Q _6081_/Y _6088_/X vssd1 vssd1 vccd1 vccd1 _6096_/Y sky130_fd_sc_hd__o21ai_1
X_9924_ _9924_/CLK _9924_/D vssd1 vssd1 vccd1 vccd1 _9924_/Q sky130_fd_sc_hd__dfxtp_1
X_5047_ _9843_/Q vssd1 vssd1 vccd1 vccd1 _5047_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9855_ _9858_/CLK _9855_/D vssd1 vssd1 vccd1 vccd1 _9855_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_198_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8806_ _8806_/A vssd1 vssd1 vccd1 vccd1 _8806_/Y sky130_fd_sc_hd__inv_2
X_9786_ _9819_/CLK _9786_/D vssd1 vssd1 vccd1 vccd1 _9786_/Q sky130_fd_sc_hd__dfxtp_1
X_6998_ _6987_/X _6997_/X _6987_/X _6997_/X vssd1 vssd1 vccd1 vccd1 _6998_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8737_ _8823_/C _8737_/B vssd1 vssd1 vccd1 vccd1 _8762_/A sky130_fd_sc_hd__or2_1
X_5949_ _9152_/X _5944_/X _9576_/Q _5945_/X vssd1 vssd1 vccd1 vccd1 _9576_/D sky130_fd_sc_hd__a22o_1
XFILLER_185_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8668_ _8668_/A vssd1 vssd1 vccd1 vccd1 _8668_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8599_ _8599_/A _8599_/B vssd1 vssd1 vccd1 vccd1 _8645_/A sky130_fd_sc_hd__or2_1
X_7619_ _7598_/A _7598_/B _7599_/B vssd1 vssd1 vccd1 vccd1 _7619_/X sky130_fd_sc_hd__a21bo_1
XFILLER_107_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7970_ _8974_/X _7987_/B vssd1 vssd1 vccd1 vccd1 _7970_/Y sky130_fd_sc_hd__nor2_1
X_6921_ _6917_/X _6918_/X _6917_/X _6918_/X vssd1 vssd1 vccd1 vccd1 _6921_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9640_ _9650_/CLK _9640_/D vssd1 vssd1 vccd1 vccd1 _9640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6852_ _6844_/X _6848_/X _6849_/X _6851_/X vssd1 vssd1 vccd1 vccd1 _6852_/X sky130_fd_sc_hd__o22a_1
X_5803_ _6567_/A _9654_/Q _5740_/Y vssd1 vssd1 vccd1 vccd1 _5803_/X sky130_fd_sc_hd__a21o_1
X_9571_ _9578_/CLK _9571_/D vssd1 vssd1 vccd1 vccd1 _9571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8522_ _8522_/A _8522_/B vssd1 vssd1 vccd1 vccd1 _8555_/A sky130_fd_sc_hd__or2_1
XFILLER_148_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6783_ _6771_/A _6771_/B _6855_/A vssd1 vssd1 vccd1 vccd1 _6786_/A sky130_fd_sc_hd__a21o_1
X_5734_ _5734_/A vssd1 vssd1 vccd1 vccd1 _8391_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8453_ _8475_/A _9377_/X vssd1 vssd1 vccd1 vccd1 _8453_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5665_ _6567_/A vssd1 vssd1 vccd1 vccd1 _8394_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_163_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8384_ _8384_/A _9679_/Q vssd1 vssd1 vccd1 vccd1 _8384_/Y sky130_fd_sc_hd__nor2_1
X_7404_ _7393_/A _7393_/B _7393_/X vssd1 vssd1 vccd1 vccd1 _7405_/B sky130_fd_sc_hd__a21bo_1
XFILLER_190_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5596_ _9706_/Q vssd1 vssd1 vccd1 vccd1 _7643_/A sky130_fd_sc_hd__inv_2
X_7335_ _9622_/Q _7408_/B _7346_/A vssd1 vssd1 vccd1 vccd1 _7336_/A sky130_fd_sc_hd__and3_1
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7266_ _7264_/X _7265_/X _7264_/X _7265_/X vssd1 vssd1 vccd1 vccd1 _7266_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_131_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9005_ _9563_/Q _9523_/Q _9013_/S vssd1 vssd1 vccd1 vccd1 _9005_/X sky130_fd_sc_hd__mux2_1
X_7197_ _7197_/A vssd1 vssd1 vccd1 vccd1 _7200_/A sky130_fd_sc_hd__inv_2
X_6217_ _8005_/A _6193_/X _6221_/C _6213_/X vssd1 vssd1 vccd1 vccd1 _6217_/Y sky130_fd_sc_hd__o22ai_1
X_6148_ _6148_/A vssd1 vssd1 vccd1 vccd1 _6148_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_12 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6079_ _7986_/A _9645_/Q _6066_/Y _6071_/A vssd1 vssd1 vccd1 vccd1 _6079_/X sky130_fd_sc_hd__o22a_1
XFILLER_57_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9907_ _9907_/CLK _9907_/D vssd1 vssd1 vccd1 vccd1 _9907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9838_ _9923_/CLK _9838_/D vssd1 vssd1 vccd1 vccd1 _9838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9769_ _9917_/CLK _9769_/D vssd1 vssd1 vccd1 vccd1 _9769_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _9907_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_177_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5450_ _7160_/A _7389_/B _6872_/A _6642_/A vssd1 vssd1 vccd1 vccd1 _5450_/X sky130_fd_sc_hd__or4_4
XFILLER_157_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5381_ _9722_/Q _5381_/B vssd1 vssd1 vccd1 vccd1 _5381_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7120_ _7120_/A _7120_/B vssd1 vssd1 vccd1 vccd1 _7121_/B sky130_fd_sc_hd__or2_1
X_7051_ _7070_/A vssd1 vssd1 vccd1 vccd1 _7051_/Y sky130_fd_sc_hd__inv_2
X_6002_ _5998_/X _6001_/X _5998_/X _6001_/X vssd1 vssd1 vccd1 vccd1 _6002_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7953_ _8807_/A vssd1 vssd1 vccd1 vccd1 _8919_/A sky130_fd_sc_hd__buf_2
XFILLER_94_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6904_ _6904_/A _6925_/B vssd1 vssd1 vccd1 vccd1 _6904_/Y sky130_fd_sc_hd__nor2_1
XPHY_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7884_ _7881_/X _7882_/B _7790_/X _7883_/Y vssd1 vssd1 vccd1 vccd1 _7884_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_35_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6835_ _6835_/A _6846_/B vssd1 vssd1 vccd1 vccd1 _6835_/Y sky130_fd_sc_hd__nor2_1
X_9623_ _9858_/CLK _9623_/D vssd1 vssd1 vccd1 vccd1 _9623_/Q sky130_fd_sc_hd__dfxtp_1
X_9554_ _9924_/CLK _9554_/D vssd1 vssd1 vccd1 vccd1 _9554_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6766_ _6766_/A _6766_/B _6766_/C vssd1 vssd1 vccd1 vccd1 _6766_/X sky130_fd_sc_hd__or3_1
XFILLER_23_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8505_ _8499_/Y _8504_/X _8499_/Y _8504_/X vssd1 vssd1 vccd1 vccd1 _8505_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_176_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5717_ _9679_/Q vssd1 vssd1 vccd1 vccd1 _5717_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6697_ _9093_/X vssd1 vssd1 vccd1 vccd1 _6764_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_9485_ _9484_/X _6978_/C _9507_/S vssd1 vssd1 vccd1 vccd1 _9485_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8436_ _9628_/Q _8580_/B _8436_/C vssd1 vssd1 vccd1 vccd1 _8436_/X sky130_fd_sc_hd__and3_1
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5648_ _9694_/Q _5645_/X _6577_/A _5635_/X _5647_/X vssd1 vssd1 vccd1 vccd1 _9694_/D
+ sky130_fd_sc_hd__o221a_1
X_8367_ _8357_/C _8366_/X _8362_/X vssd1 vssd1 vccd1 vccd1 _8367_/X sky130_fd_sc_hd__o21a_1
X_5579_ _5579_/A _5579_/B vssd1 vssd1 vccd1 vccd1 _9710_/D sky130_fd_sc_hd__nor2_1
X_8298_ _4770_/X _8198_/X _8297_/X vssd1 vssd1 vccd1 vccd1 _8298_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_144_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7318_ _9475_/X vssd1 vssd1 vccd1 vccd1 _7321_/B sky130_fd_sc_hd__inv_2
XFILLER_131_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7249_ _7249_/A vssd1 vssd1 vccd1 vccd1 _7249_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput8 io_wb_adr_i[3] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_4
XFILLER_64_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4950_ _9117_/X _4943_/X _9854_/Q _4944_/X _4947_/X vssd1 vssd1 vccd1 vccd1 _9854_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_205_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4881_ _5206_/A vssd1 vssd1 vccd1 vccd1 _4881_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_189_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6620_ _6620_/A vssd1 vssd1 vccd1 vccd1 _6691_/C sky130_fd_sc_hd__inv_2
XFILLER_32_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6551_ _6558_/A vssd1 vssd1 vccd1 vccd1 _6551_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5502_ _9383_/X _5501_/X _9383_/X _5501_/X vssd1 vssd1 vccd1 vccd1 _5605_/A sky130_fd_sc_hd__a2bb2oi_1
X_6482_ _6368_/X _6481_/X _6368_/X _6481_/X vssd1 vssd1 vccd1 vccd1 _6482_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_118_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9270_ _9269_/X input18/X _9282_/S vssd1 vssd1 vccd1 vccd1 _9270_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8221_ _8221_/A _8227_/B vssd1 vssd1 vccd1 vccd1 _8221_/X sky130_fd_sc_hd__or2_1
X_5433_ _9345_/X vssd1 vssd1 vccd1 vccd1 _5434_/B sky130_fd_sc_hd__inv_2
XFILLER_145_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8152_ _7713_/X _8113_/Y _7840_/A _8110_/X _8151_/X vssd1 vssd1 vccd1 vccd1 _8152_/X
+ sky130_fd_sc_hd__o221a_1
X_5364_ _5364_/A vssd1 vssd1 vccd1 vccd1 _5364_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7103_ _9620_/Q vssd1 vssd1 vccd1 vccd1 _7324_/A sky130_fd_sc_hd__inv_2
XFILLER_206_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8083_ _9555_/Q _8083_/B vssd1 vssd1 vccd1 vccd1 _8084_/B sky130_fd_sc_hd__or2_2
XFILLER_141_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5295_ _9737_/Q _5295_/B vssd1 vssd1 vccd1 vccd1 _5295_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7034_ _7016_/X _7017_/X _7018_/X _7033_/X vssd1 vssd1 vccd1 vccd1 _7034_/X sky130_fd_sc_hd__o22a_1
XFILLER_142_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8985_ _6453_/A _7755_/X _9480_/S vssd1 vssd1 vccd1 vccd1 _8985_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7936_ _9494_/X _7956_/B vssd1 vssd1 vccd1 vccd1 _7936_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7867_ _7865_/A _7865_/B _7839_/X _7866_/Y vssd1 vssd1 vccd1 vccd1 _7867_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_35_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6818_ _6806_/A _6806_/B _6806_/X vssd1 vssd1 vccd1 vccd1 _6819_/B sky130_fd_sc_hd__a21bo_1
XPHY_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9606_ _9895_/CLK _9606_/D vssd1 vssd1 vccd1 vccd1 _9606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7798_ _7803_/B vssd1 vssd1 vccd1 vccd1 _7798_/Y sky130_fd_sc_hd__inv_2
XPHY_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9537_ _9907_/CLK _9537_/D vssd1 vssd1 vccd1 vccd1 _9537_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6749_ _6749_/A _6748_/X vssd1 vssd1 vccd1 vccd1 _6749_/X sky130_fd_sc_hd__or2b_1
XFILLER_183_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9468_ _7038_/Y _7082_/Y _9683_/Q vssd1 vssd1 vccd1 vccd1 _9468_/X sky130_fd_sc_hd__mux2_1
X_8419_ _8543_/B _8415_/X _8432_/B vssd1 vssd1 vccd1 vccd1 _8419_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_191_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9399_ _8003_/X _6101_/Y _9504_/S vssd1 vssd1 vccd1 vccd1 _9399_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5080_ _9804_/Q vssd1 vssd1 vccd1 vccd1 _6317_/D sky130_fd_sc_hd__inv_2
XFILLER_96_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_34_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _9895_/CLK sky130_fd_sc_hd__clkbuf_16
X_8770_ _8942_/A _8893_/B _8609_/A _8769_/X vssd1 vssd1 vccd1 vccd1 _8770_/X sky130_fd_sc_hd__o31a_1
X_5982_ _5701_/A _9635_/Q _5981_/A _5704_/B _5981_/Y vssd1 vssd1 vccd1 vccd1 _5982_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_64_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7721_ _9914_/Q vssd1 vssd1 vccd1 vccd1 _7848_/A sky130_fd_sc_hd__inv_2
XFILLER_17_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4933_ _4952_/A vssd1 vssd1 vccd1 vccd1 _4951_/A sky130_fd_sc_hd__inv_2
XFILLER_205_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7652_ _7652_/A _7652_/B vssd1 vssd1 vccd1 vccd1 _7652_/Y sky130_fd_sc_hd__nor2_1
X_4864_ _4880_/A vssd1 vssd1 vccd1 vccd1 _4879_/A sky130_fd_sc_hd__inv_2
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4795_ _9302_/X _4782_/X _4794_/X _4784_/X _4791_/X vssd1 vssd1 vccd1 vccd1 _9919_/D
+ sky130_fd_sc_hd__o221a_1
X_6603_ _6730_/A vssd1 vssd1 vccd1 vccd1 _6971_/A sky130_fd_sc_hd__buf_2
X_7583_ _7583_/A vssd1 vssd1 vccd1 vccd1 _7599_/A sky130_fd_sc_hd__inv_2
X_9322_ _9321_/X input36/X _9334_/S vssd1 vssd1 vccd1 vccd1 _9322_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6534_ _6535_/A _6534_/B vssd1 vssd1 vccd1 vccd1 _6534_/Y sky130_fd_sc_hd__nor2_1
XFILLER_192_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9253_ _9252_/X _7808_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9253_/X sky130_fd_sc_hd__mux2_1
X_6465_ _6432_/Y _6465_/B _6465_/C _6465_/D vssd1 vssd1 vccd1 vccd1 _6466_/D sky130_fd_sc_hd__and4b_1
XFILLER_173_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8204_ _8204_/A _8204_/B vssd1 vssd1 vccd1 vccd1 _8205_/B sky130_fd_sc_hd__nand2_1
XFILLER_161_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5416_ _9363_/X vssd1 vssd1 vccd1 vccd1 _5418_/A sky130_fd_sc_hd__inv_2
X_6396_ _9778_/Q _8197_/A vssd1 vssd1 vccd1 vccd1 _6397_/A sky130_fd_sc_hd__or2_2
XFILLER_161_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9184_ _6525_/Y _9789_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9538_/D sky130_fd_sc_hd__mux2_1
X_8135_ _8133_/X _8134_/Y _7657_/A _8126_/Y vssd1 vssd1 vccd1 vccd1 _8135_/X sky130_fd_sc_hd__o22a_1
XFILLER_121_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5347_ _9729_/Q _5347_/B vssd1 vssd1 vccd1 vccd1 _5347_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8066_ _9538_/Q _8066_/B vssd1 vssd1 vccd1 vccd1 _8067_/B sky130_fd_sc_hd__or2_1
XFILLER_99_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5278_ _5278_/A vssd1 vssd1 vccd1 vccd1 _5279_/B sky130_fd_sc_hd__inv_2
X_7017_ _6620_/A _7001_/X _6620_/A _7001_/X vssd1 vssd1 vccd1 vccd1 _7017_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8968_ _4753_/A _8967_/X _9930_/Q _4753_/Y _5891_/X vssd1 vssd1 vccd1 vccd1 _9930_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_83_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7919_ _7919_/A vssd1 vssd1 vccd1 vccd1 _8046_/B sky130_fd_sc_hd__buf_4
XFILLER_196_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8899_ _8859_/X _8898_/X _8859_/X _8898_/X vssd1 vssd1 vccd1 vccd1 _8899_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput22 io_wb_dat_i[15] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_6
Xinput11 io_wb_adr_i[6] vssd1 vssd1 vccd1 vccd1 _5707_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_190_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput33 io_wb_dat_i[25] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_4
XPHY_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput44 io_wb_dat_i[6] vssd1 vssd1 vccd1 vccd1 _5029_/A sky130_fd_sc_hd__buf_4
XFILLER_155_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6250_ _9584_/Q vssd1 vssd1 vccd1 vccd1 _8024_/A sky130_fd_sc_hd__inv_2
XFILLER_115_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5201_ input17/X _5192_/X _6337_/A _5193_/X _5194_/X vssd1 vssd1 vccd1 vccd1 _9758_/D
+ sky130_fd_sc_hd__a221o_1
X_6181_ _9572_/Q vssd1 vssd1 vccd1 vccd1 _7983_/A sky130_fd_sc_hd__inv_2
X_5132_ _5165_/A vssd1 vssd1 vccd1 vccd1 _5132_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5063_ _9840_/Q vssd1 vssd1 vccd1 vccd1 _5063_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9871_ _9893_/CLK _9871_/D vssd1 vssd1 vccd1 vccd1 _9871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8822_ _8865_/C vssd1 vssd1 vccd1 vccd1 _8901_/C sky130_fd_sc_hd__inv_2
XFILLER_92_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8753_ _9395_/X vssd1 vssd1 vccd1 vccd1 _8821_/B sky130_fd_sc_hd__clkbuf_2
X_5965_ _9142_/X _5937_/A _9564_/Q _5938_/A vssd1 vssd1 vccd1 vccd1 _9564_/D sky130_fd_sc_hd__a22o_1
XFILLER_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8684_ _9439_/X vssd1 vssd1 vccd1 vccd1 _8751_/B sky130_fd_sc_hd__clkbuf_2
X_7704_ _4820_/X _6335_/Y _7861_/A _6350_/A _7703_/X vssd1 vssd1 vccd1 vccd1 _7705_/D
+ sky130_fd_sc_hd__o221a_1
X_5896_ _6756_/A _5884_/A _5039_/A _5885_/A _5891_/X vssd1 vssd1 vccd1 vccd1 _9612_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_80_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4916_ _9871_/Q _4914_/X _9723_/Q _4912_/X _4915_/X vssd1 vssd1 vccd1 vccd1 _9871_/D
+ sky130_fd_sc_hd__o221a_1
X_4847_ _9899_/Q vssd1 vssd1 vccd1 vccd1 _4847_/X sky130_fd_sc_hd__clkbuf_2
X_7635_ _7644_/A vssd1 vssd1 vccd1 vccd1 _7640_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_138_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9305_ _9304_/X _7878_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9305_/X sky130_fd_sc_hd__mux2_1
X_4778_ _4830_/A vssd1 vssd1 vccd1 vccd1 _4778_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_153_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7566_ _7542_/X _7549_/X _7542_/X _7549_/X vssd1 vssd1 vccd1 vccd1 _7582_/A sky130_fd_sc_hd__a2bb2o_1
X_6517_ _6316_/B _6401_/Y _6316_/A _6399_/Y _6516_/X vssd1 vssd1 vccd1 vccd1 _6517_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7497_ _7497_/A _9432_/X vssd1 vssd1 vccd1 vccd1 _7497_/X sky130_fd_sc_hd__or2_1
X_9236_ _9751_/Q _9235_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9236_/X sky130_fd_sc_hd__mux2_1
X_6448_ _9789_/Q _6525_/B vssd1 vssd1 vccd1 vccd1 _6448_/Y sky130_fd_sc_hd__nor2_1
X_9167_ _6289_/Y input36/X _9170_/S vssd1 vssd1 vccd1 vccd1 _9167_/X sky130_fd_sc_hd__mux2_1
X_6379_ _9761_/Q _6435_/A vssd1 vssd1 vccd1 vccd1 _8229_/A sky130_fd_sc_hd__or2_2
X_8118_ _9538_/Q _8066_/B _8067_/B vssd1 vssd1 vccd1 vccd1 _8118_/X sky130_fd_sc_hd__a21bo_1
XFILLER_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9098_ _6000_/X _6002_/X _9896_/Q vssd1 vssd1 vccd1 vccd1 _9098_/X sky130_fd_sc_hd__mux2_1
X_8049_ _9533_/Q vssd1 vssd1 vccd1 vccd1 _8324_/B sky130_fd_sc_hd__inv_2
XFILLER_87_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5750_ _6558_/A _9658_/Q _5731_/Y _5749_/X vssd1 vssd1 vccd1 vccd1 _5750_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5681_ _5689_/A vssd1 vssd1 vccd1 vccd1 _5681_/X sky130_fd_sc_hd__buf_1
XFILLER_30_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7420_ _7420_/A _7420_/B vssd1 vssd1 vccd1 vccd1 _7442_/B sky130_fd_sc_hd__nor2_2
XFILLER_190_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7351_ _7351_/A vssd1 vssd1 vccd1 vccd1 _7352_/A sky130_fd_sc_hd__inv_2
X_6302_ _6171_/X _6301_/X _6171_/X _6301_/X vssd1 vssd1 vccd1 vccd1 _6302_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_190_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7282_ _7282_/A vssd1 vssd1 vccd1 vccd1 _7283_/C sky130_fd_sc_hd__inv_2
XFILLER_170_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9021_ _9785_/Q _9902_/Q _9480_/S vssd1 vssd1 vccd1 vccd1 _9021_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6233_ _8013_/A _6139_/A _8015_/A _6139_/A vssd1 vssd1 vccd1 vccd1 _6234_/B sky130_fd_sc_hd__o22a_1
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6164_ _9570_/Q _6165_/A _7973_/A _6148_/X vssd1 vssd1 vccd1 vccd1 _6176_/A sky130_fd_sc_hd__a22o_1
X_5115_ _5115_/A _5115_/B vssd1 vssd1 vccd1 vccd1 _9797_/D sky130_fd_sc_hd__nor2_1
XFILLER_97_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6095_ _6095_/A _6095_/B vssd1 vssd1 vccd1 vccd1 _6095_/X sky130_fd_sc_hd__or2_1
XFILLER_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5046_ _9811_/Q vssd1 vssd1 vccd1 vccd1 _6316_/A sky130_fd_sc_hd__inv_2
X_9923_ _9923_/CLK _9923_/D vssd1 vssd1 vccd1 vccd1 _9923_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9854_ _9858_/CLK _9854_/D vssd1 vssd1 vccd1 vccd1 _9854_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8805_ _8805_/A _8778_/X vssd1 vssd1 vccd1 vccd1 _8806_/A sky130_fd_sc_hd__or2b_1
X_9785_ _9819_/CLK _9785_/D vssd1 vssd1 vccd1 vccd1 _9785_/Q sky130_fd_sc_hd__dfxtp_1
X_6997_ _6989_/X _6993_/X _6995_/X _6996_/X vssd1 vssd1 vccd1 vccd1 _6997_/X sky130_fd_sc_hd__o22a_1
XFILLER_53_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8736_ _8734_/X _8735_/X _8734_/X _8735_/X vssd1 vssd1 vccd1 vccd1 _8737_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5948_ _9153_/X _5944_/X _9577_/Q _5945_/X vssd1 vssd1 vccd1 vccd1 _9577_/D sky130_fd_sc_hd__a22o_1
XFILLER_178_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8667_ _8665_/Y _8666_/Y _8665_/Y _8666_/Y vssd1 vssd1 vccd1 vccd1 _8667_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_166_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5879_ _9619_/Q vssd1 vssd1 vccd1 vccd1 _7492_/C sky130_fd_sc_hd__buf_2
XFILLER_154_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8598_ _8599_/B vssd1 vssd1 vccd1 vccd1 _8598_/Y sky130_fd_sc_hd__inv_2
X_7618_ _7075_/A _7075_/B _7076_/B vssd1 vssd1 vccd1 vccd1 _7618_/X sky130_fd_sc_hd__a21bo_1
XFILLER_153_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7549_ _7543_/X _7545_/X _7546_/X _7548_/X vssd1 vssd1 vccd1 vccd1 _7549_/X sky130_fd_sc_hd__o22a_1
XFILLER_153_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9219_ _9824_/Q _7650_/Y _9528_/Q vssd1 vssd1 vccd1 vccd1 _9219_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6920_ _6914_/X _6919_/X _6914_/X _6919_/X vssd1 vssd1 vccd1 vccd1 _6920_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_207_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6851_ _6851_/A _6851_/B vssd1 vssd1 vccd1 vccd1 _6851_/X sky130_fd_sc_hd__or2_1
X_5802_ _9655_/Q _5793_/X _5787_/X _7086_/A _5791_/X vssd1 vssd1 vccd1 vccd1 _9655_/D
+ sky130_fd_sc_hd__o221a_1
X_9570_ _9578_/CLK _9570_/D vssd1 vssd1 vccd1 vccd1 _9570_/Q sky130_fd_sc_hd__dfxtp_1
X_8521_ _8521_/A vssd1 vssd1 vccd1 vccd1 _8522_/B sky130_fd_sc_hd__inv_2
X_6782_ _6782_/A vssd1 vssd1 vccd1 vccd1 _6855_/A sky130_fd_sc_hd__inv_2
XFILLER_148_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5733_ _9673_/Q vssd1 vssd1 vccd1 vccd1 _5734_/A sky130_fd_sc_hd__inv_2
X_8452_ _8452_/A _9378_/X vssd1 vssd1 vccd1 vccd1 _8452_/X sky130_fd_sc_hd__or2_1
XFILLER_175_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5664_ _9671_/Q vssd1 vssd1 vccd1 vccd1 _6567_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5595_ _5595_/A _5595_/B vssd1 vssd1 vccd1 vccd1 _5595_/Y sky130_fd_sc_hd__nor2_1
X_8383_ _9695_/Q vssd1 vssd1 vccd1 vccd1 _8384_/A sky130_fd_sc_hd__inv_2
X_7403_ _7403_/A _7384_/X vssd1 vssd1 vccd1 vccd1 _7405_/A sky130_fd_sc_hd__or2b_1
XFILLER_163_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7334_ _7334_/A _7334_/B vssd1 vssd1 vccd1 vccd1 _7346_/A sky130_fd_sc_hd__or2_1
XFILLER_131_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7265_ _7265_/A _9470_/X vssd1 vssd1 vccd1 vccd1 _7265_/X sky130_fd_sc_hd__or2_1
X_9004_ _9003_/X _9748_/Q _9481_/S vssd1 vssd1 vccd1 vccd1 _9004_/X sky130_fd_sc_hd__mux2_2
XFILLER_131_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7196_ _7497_/A _9414_/X _7201_/A _9415_/X vssd1 vssd1 vccd1 vccd1 _7197_/A sky130_fd_sc_hd__or4_4
X_6216_ _9578_/Q _6166_/A _8010_/A _6201_/A vssd1 vssd1 vccd1 vccd1 _6221_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6147_ _9567_/Q vssd1 vssd1 vccd1 vccd1 _7949_/A sky130_fd_sc_hd__inv_2
XINSDIODE2_13 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6078_ _6076_/Y _6077_/X _6076_/Y _6077_/X vssd1 vssd1 vccd1 vccd1 _6078_/X sky130_fd_sc_hd__a2bb2o_1
X_9906_ _9917_/CLK _9906_/D vssd1 vssd1 vccd1 vccd1 _9906_/Q sky130_fd_sc_hd__dfxtp_2
X_5029_ _5029_/A vssd1 vssd1 vccd1 vccd1 _5029_/X sky130_fd_sc_hd__buf_4
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9837_ _9923_/CLK _9837_/D vssd1 vssd1 vccd1 vccd1 _9837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9768_ _9917_/CLK _9768_/D vssd1 vssd1 vccd1 vccd1 _9768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8719_ _8710_/X _8718_/X _8710_/X _8718_/X vssd1 vssd1 vccd1 vccd1 _8719_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_139_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9699_ _9699_/CLK _9699_/D vssd1 vssd1 vccd1 vccd1 _9699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5380_ _5380_/A vssd1 vssd1 vccd1 vccd1 _5381_/B sky130_fd_sc_hd__inv_2
XFILLER_153_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7050_ _6834_/A _6834_/B _6846_/B vssd1 vssd1 vccd1 vccd1 _7070_/A sky130_fd_sc_hd__a21oi_2
XFILLER_101_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6001_ _7935_/A _9637_/Q _5989_/A _5992_/A vssd1 vssd1 vccd1 vccd1 _6001_/X sky130_fd_sc_hd__o22a_1
XFILLER_39_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7952_ _8776_/A vssd1 vssd1 vccd1 vccd1 _8807_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6903_ _6903_/A _6903_/B vssd1 vssd1 vccd1 vccd1 _6925_/B sky130_fd_sc_hd__nor2_2
XFILLER_211_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7883_ _7887_/B vssd1 vssd1 vccd1 vccd1 _7883_/Y sky130_fd_sc_hd__inv_2
X_9622_ _9715_/CLK _9622_/D vssd1 vssd1 vccd1 vccd1 _9622_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_211_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6834_ _6834_/A _6834_/B vssd1 vssd1 vccd1 vccd1 _6846_/B sky130_fd_sc_hd__nor2_2
XFILLER_62_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9553_ _9924_/CLK _9553_/D vssd1 vssd1 vccd1 vccd1 _9553_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6765_ _6765_/A vssd1 vssd1 vccd1 vccd1 _6766_/C sky130_fd_sc_hd__inv_2
XFILLER_23_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8504_ _8823_/A _8500_/Y _8529_/C _8503_/X vssd1 vssd1 vccd1 vccd1 _8504_/X sky130_fd_sc_hd__a31o_1
X_5716_ _9680_/Q _9663_/Q vssd1 vssd1 vccd1 vccd1 _5716_/Y sky130_fd_sc_hd__nor2_1
X_9484_ _9483_/X _7518_/A _9506_/S vssd1 vssd1 vccd1 vccd1 _9484_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8435_ _8452_/A _9377_/X vssd1 vssd1 vccd1 vccd1 _8475_/C sky130_fd_sc_hd__nor2_4
XFILLER_176_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6696_ _6883_/A vssd1 vssd1 vccd1 vccd1 _7005_/A sky130_fd_sc_hd__buf_4
XFILLER_191_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5647_ _5660_/A vssd1 vssd1 vccd1 vccd1 _5647_/X sky130_fd_sc_hd__clkbuf_2
X_8366_ _4780_/X _8359_/Y _4775_/X _8354_/Y _8365_/Y vssd1 vssd1 vccd1 vccd1 _8366_/X
+ sky130_fd_sc_hd__o221a_1
X_5578_ _5553_/X _5573_/Y _5574_/Y _7648_/A _5577_/X vssd1 vssd1 vccd1 vccd1 _5579_/B
+ sky130_fd_sc_hd__o32a_1
X_8297_ _7902_/A _8201_/Y _8296_/X vssd1 vssd1 vccd1 vccd1 _8297_/X sky130_fd_sc_hd__a21o_1
XFILLER_151_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7317_ _7317_/A _7379_/A vssd1 vssd1 vccd1 vccd1 _7324_/C sky130_fd_sc_hd__nor2_2
X_7248_ _9626_/Q _7291_/B _7259_/A vssd1 vssd1 vccd1 vccd1 _7249_/A sky130_fd_sc_hd__and3_1
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7179_ _9622_/Q _7210_/B _7190_/A vssd1 vssd1 vccd1 vccd1 _7180_/A sky130_fd_sc_hd__and3_1
XFILLER_58_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 io_wb_adr_i[4] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_1
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4880_ _4880_/A vssd1 vssd1 vccd1 vccd1 _4880_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6550_ _6550_/A _6550_/B vssd1 vssd1 vccd1 vccd1 _6550_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5501_ _5428_/X _5453_/X _5428_/X _5453_/X vssd1 vssd1 vccd1 vccd1 _5501_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_173_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6481_ _8184_/A _8183_/B _6363_/Y vssd1 vssd1 vccd1 vccd1 _6481_/X sky130_fd_sc_hd__a21o_1
XFILLER_145_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8220_ _5181_/X _8219_/X _8216_/B vssd1 vssd1 vccd1 vccd1 _8220_/X sky130_fd_sc_hd__a21bo_1
X_5432_ _9347_/X vssd1 vssd1 vccd1 vccd1 _5434_/A sky130_fd_sc_hd__inv_2
XFILLER_160_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8151_ _7835_/A _8113_/Y _7698_/X _8114_/X _8150_/X vssd1 vssd1 vccd1 vccd1 _8151_/X
+ sky130_fd_sc_hd__a221o_1
X_5363_ _5363_/A vssd1 vssd1 vccd1 vccd1 _5364_/A sky130_fd_sc_hd__clkbuf_2
X_7102_ _7101_/X _5811_/Y _7084_/B vssd1 vssd1 vccd1 vccd1 _7102_/Y sky130_fd_sc_hd__o21ai_1
X_8082_ _9554_/Q _8082_/B vssd1 vssd1 vccd1 vccd1 _8083_/B sky130_fd_sc_hd__or2_1
XFILLER_113_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5294_ _5294_/A vssd1 vssd1 vccd1 vccd1 _5295_/B sky130_fd_sc_hd__inv_2
XFILLER_141_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7033_ _7019_/X _7020_/X _7021_/X _7032_/X vssd1 vssd1 vccd1 vccd1 _7033_/X sky130_fd_sc_hd__o22a_1
XFILLER_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8984_ _8983_/X _7005_/A _9507_/S vssd1 vssd1 vccd1 vccd1 _8984_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7935_ _7935_/A _9503_/S vssd1 vssd1 vccd1 vccd1 _7935_/X sky130_fd_sc_hd__or2_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7866_ _7869_/B vssd1 vssd1 vccd1 vccd1 _7866_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6817_ _6817_/A _6796_/X vssd1 vssd1 vccd1 vccd1 _6819_/A sky130_fd_sc_hd__or2b_1
XPHY_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9605_ _9895_/CLK _9605_/D vssd1 vssd1 vccd1 vccd1 _9605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7797_ _7797_/A _7797_/B vssd1 vssd1 vccd1 vccd1 _7803_/B sky130_fd_sc_hd__or2_1
X_9536_ _9796_/CLK _9536_/D vssd1 vssd1 vccd1 vccd1 _9536_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6748_ _6764_/A _6760_/B _6766_/A _6764_/B vssd1 vssd1 vccd1 vccd1 _6748_/X sky130_fd_sc_hd__or4_4
XFILLER_176_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9467_ _6598_/X _6599_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9467_/X sky130_fd_sc_hd__mux2_2
X_6679_ _6978_/A vssd1 vssd1 vccd1 vccd1 _6982_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_191_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8418_ _5515_/X _6890_/A _8397_/Y vssd1 vssd1 vccd1 vccd1 _8432_/B sky130_fd_sc_hd__o21ai_4
XFILLER_109_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9398_ _9397_/X _9763_/Q _9481_/S vssd1 vssd1 vccd1 vccd1 _9398_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8349_ _7673_/A _8342_/Y _4802_/X _8337_/Y _8348_/Y vssd1 vssd1 vccd1 vccd1 _8349_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_117_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_0_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _9909_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5981_ _5981_/A vssd1 vssd1 vccd1 vccd1 _5981_/Y sky130_fd_sc_hd__inv_2
X_7720_ _7769_/A _6341_/Y _7887_/A _8205_/A _7719_/X vssd1 vssd1 vccd1 vccd1 _7731_/C
+ sky130_fd_sc_hd__o221a_1
X_4932_ _5816_/A _5967_/A _9667_/Q vssd1 vssd1 vccd1 vccd1 _4952_/A sky130_fd_sc_hd__o21ai_4
XFILLER_205_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7651_ _7651_/A _7652_/B vssd1 vssd1 vccd1 vccd1 _7651_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6602_ _6890_/B vssd1 vssd1 vccd1 vccd1 _6730_/A sky130_fd_sc_hd__buf_1
X_4863_ _5222_/A _9335_/X vssd1 vssd1 vccd1 vccd1 _4880_/A sky130_fd_sc_hd__or2_4
XFILLER_32_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4794_ _4794_/A vssd1 vssd1 vccd1 vccd1 _4794_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7582_ _7582_/A vssd1 vssd1 vccd1 vccd1 _7600_/A sky130_fd_sc_hd__inv_2
XFILLER_32_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9321_ _9320_/X _7898_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9321_/X sky130_fd_sc_hd__mux2_1
X_6533_ _6535_/A _6533_/B vssd1 vssd1 vccd1 vccd1 _6533_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9252_ _9755_/Q _9251_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9252_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6464_ _9795_/Q _6532_/B vssd1 vssd1 vccd1 vccd1 _6465_/D sky130_fd_sc_hd__nand2_1
XFILLER_173_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8203_ _8203_/A _8211_/B vssd1 vssd1 vccd1 vccd1 _8204_/B sky130_fd_sc_hd__nor2_1
X_5415_ _5415_/A _5415_/B vssd1 vssd1 vccd1 vccd1 _5415_/Y sky130_fd_sc_hd__nor2_1
X_6395_ _9777_/Q _6402_/A vssd1 vssd1 vccd1 vccd1 _8197_/A sky130_fd_sc_hd__or2_2
XFILLER_161_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9183_ _6522_/Y _9788_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9537_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8134_ _8134_/A _8134_/B vssd1 vssd1 vccd1 vccd1 _8134_/Y sky130_fd_sc_hd__nor2_1
X_5346_ _5346_/A vssd1 vssd1 vccd1 vccd1 _5347_/B sky130_fd_sc_hd__inv_2
X_8065_ _9537_/Q _8065_/B vssd1 vssd1 vccd1 vccd1 _8066_/B sky130_fd_sc_hd__or2_2
XFILLER_102_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5277_ _5277_/A vssd1 vssd1 vccd1 vccd1 _9742_/D sky130_fd_sc_hd__inv_2
X_7016_ _6913_/X _6960_/X _6913_/X _6960_/X vssd1 vssd1 vccd1 vccd1 _7016_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8967_ _9527_/Q _8967_/B vssd1 vssd1 vccd1 vccd1 _8967_/X sky130_fd_sc_hd__and2_1
XFILLER_16_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7918_ _7918_/A _7918_/B vssd1 vssd1 vccd1 vccd1 _9051_/S sky130_fd_sc_hd__nor2_8
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8898_ _8894_/Y _8897_/Y _8894_/Y _8897_/Y vssd1 vssd1 vccd1 vccd1 _8898_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_70_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7849_ _7852_/B vssd1 vssd1 vccd1 vccd1 _7849_/Y sky130_fd_sc_hd__inv_2
XPHY_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9519_ _9519_/CLK input2/X vssd1 vssd1 vccd1 vccd1 _9520_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput12 io_wb_adr_i[7] vssd1 vssd1 vccd1 vccd1 _5707_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_190_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput34 io_wb_dat_i[26] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_4
Xinput23 io_wb_dat_i[16] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_4
XPHY_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput45 io_wb_dat_i[7] vssd1 vssd1 vccd1 vccd1 _5026_/A sky130_fd_sc_hd__buf_6
XFILLER_170_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5200_ _9758_/Q vssd1 vssd1 vccd1 vccd1 _6337_/A sky130_fd_sc_hd__buf_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6180_ _6179_/A _6179_/B _6187_/A vssd1 vssd1 vccd1 vccd1 _6180_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_130_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5131_ _5128_/X _9790_/Q _5130_/X _9217_/X _5124_/X vssd1 vssd1 vccd1 vccd1 _9790_/D
+ sky130_fd_sc_hd__o221a_1
X_5062_ _9808_/Q vssd1 vssd1 vccd1 vccd1 _6316_/D sky130_fd_sc_hd__inv_2
XFILLER_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9870_ _9893_/CLK _9870_/D vssd1 vssd1 vccd1 vccd1 _9870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8821_ _8821_/A _8821_/B vssd1 vssd1 vccd1 vccd1 _8865_/C sky130_fd_sc_hd__or2_2
XFILLER_65_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8752_ _8752_/A _8751_/X vssd1 vssd1 vccd1 vccd1 _8760_/A sky130_fd_sc_hd__or2b_1
XFILLER_80_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7703_ _9915_/Q _6351_/Y _4765_/A _6354_/Y vssd1 vssd1 vccd1 vccd1 _7703_/X sky130_fd_sc_hd__o22a_1
X_5964_ _9075_/X _5958_/X _9565_/Q _5959_/X vssd1 vssd1 vccd1 vccd1 _9565_/D sky130_fd_sc_hd__a22o_1
X_8683_ _8640_/Y _8682_/X _8640_/Y _8682_/X vssd1 vssd1 vccd1 vccd1 _8683_/X sky130_fd_sc_hd__a2bb2o_1
X_5895_ _9612_/Q vssd1 vssd1 vccd1 vccd1 _6756_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4915_ _4923_/A vssd1 vssd1 vccd1 vccd1 _4915_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4846_ _9238_/X _4834_/X _4843_/X _4836_/X _4845_/X vssd1 vssd1 vccd1 vccd1 _9900_/D
+ sky130_fd_sc_hd__o221a_1
X_7634_ _9715_/Q _9350_/X vssd1 vssd1 vccd1 vccd1 _7644_/A sky130_fd_sc_hd__or2b_2
XFILLER_178_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7565_ _7539_/X _7550_/X _7539_/X _7550_/X vssd1 vssd1 vccd1 vccd1 _7581_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6516_ _6316_/B _6401_/Y _6316_/C _6405_/A _6515_/Y vssd1 vssd1 vccd1 vccd1 _6516_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_165_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9304_ _9772_/Q _9303_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9304_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4777_ _5405_/A vssd1 vssd1 vccd1 vccd1 _4830_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_180_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7496_ _7490_/X _7495_/X _7490_/X _7495_/X vssd1 vssd1 vccd1 vccd1 _7496_/X sky130_fd_sc_hd__a2bb2o_1
X_9235_ _7787_/X _9751_/Q _9327_/S vssd1 vssd1 vccd1 vccd1 _9235_/X sky130_fd_sc_hd__mux2_1
X_6447_ _6447_/A vssd1 vssd1 vccd1 vccd1 _6525_/B sky130_fd_sc_hd__inv_2
X_9166_ _6282_/X input35/X _9170_/S vssd1 vssd1 vccd1 vccd1 _9166_/X sky130_fd_sc_hd__mux2_1
X_6378_ _9760_/Q _8231_/A vssd1 vssd1 vccd1 vccd1 _6435_/A sky130_fd_sc_hd__or2_1
XFILLER_88_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8117_ _9539_/Q _8067_/B _8068_/B vssd1 vssd1 vccd1 vccd1 _8117_/X sky130_fd_sc_hd__a21bo_1
X_5329_ _5329_/A _5380_/A vssd1 vssd1 vccd1 vccd1 _5375_/A sky130_fd_sc_hd__or2_1
XFILLER_87_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9097_ _5990_/Y _5993_/X _9896_/Q vssd1 vssd1 vccd1 vccd1 _9097_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8048_ _9559_/Q vssd1 vssd1 vccd1 vccd1 _8048_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_33_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _9888_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5680_ _6596_/A _5671_/X _9107_/X _5676_/X _5674_/X vssd1 vssd1 vccd1 vccd1 _9680_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_175_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7350_ _7350_/A _7350_/B vssd1 vssd1 vccd1 vccd1 _7350_/X sky130_fd_sc_hd__or2_1
X_6301_ _8046_/A _6300_/X _8046_/A _6300_/X vssd1 vssd1 vccd1 vccd1 _6301_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_128_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7281_ _7290_/A _9470_/X vssd1 vssd1 vccd1 vccd1 _7282_/A sky130_fd_sc_hd__or2_2
X_6232_ _6232_/A _6232_/B vssd1 vssd1 vccd1 vccd1 _6244_/C sky130_fd_sc_hd__or2_1
X_9020_ _7949_/Y _9599_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9020_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6163_ _9570_/Q vssd1 vssd1 vccd1 vccd1 _7973_/A sky130_fd_sc_hd__inv_2
X_5114_ _5128_/A _5112_/Y _5113_/Y _5097_/X vssd1 vssd1 vccd1 vccd1 _5115_/B sky130_fd_sc_hd__o22a_1
X_6094_ _9861_/Q _6094_/B vssd1 vssd1 vccd1 vccd1 _6095_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9922_ _9923_/CLK _9922_/D vssd1 vssd1 vccd1 vccd1 _9922_/Q sky130_fd_sc_hd__dfxtp_1
X_5045_ _5136_/A vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__buf_2
XFILLER_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9853_ _9879_/CLK _9853_/D vssd1 vssd1 vccd1 vccd1 _9853_/Q sky130_fd_sc_hd__dfxtp_2
X_8804_ _8893_/C _8803_/A _8801_/A _8803_/Y vssd1 vssd1 vccd1 vccd1 _8804_/X sky130_fd_sc_hd__a22o_2
X_9784_ _9819_/CLK _9784_/D vssd1 vssd1 vccd1 vccd1 _9784_/Q sky130_fd_sc_hd__dfxtp_1
X_6996_ _6989_/X _6993_/X _6989_/X _6993_/X vssd1 vssd1 vccd1 vccd1 _6996_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_198_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8735_ _8735_/A _9439_/X _8735_/C vssd1 vssd1 vccd1 vccd1 _8735_/X sky130_fd_sc_hd__or3_1
XFILLER_80_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5947_ _9154_/X _5944_/X _9578_/Q _5945_/X vssd1 vssd1 vccd1 vccd1 _9578_/D sky130_fd_sc_hd__a22o_1
X_8666_ _8621_/A _8620_/Y _8709_/A vssd1 vssd1 vccd1 vccd1 _8666_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5878_ _7273_/A _5865_/A _5039_/X _5866_/A _5875_/X vssd1 vssd1 vccd1 vccd1 _9620_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7617_ _7599_/A _7599_/B _7600_/B vssd1 vssd1 vccd1 vccd1 _7617_/X sky130_fd_sc_hd__a21bo_1
X_8597_ _8596_/A _8596_/B _8596_/Y vssd1 vssd1 vccd1 vccd1 _8599_/B sky130_fd_sc_hd__a21oi_4
XFILLER_166_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4829_ _7810_/A vssd1 vssd1 vccd1 vccd1 _7769_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7548_ _7548_/A _7548_/B vssd1 vssd1 vccd1 vccd1 _7548_/X sky130_fd_sc_hd__or2_1
XFILLER_134_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7479_ _7426_/X _7429_/X _7430_/X _7478_/X vssd1 vssd1 vccd1 vccd1 _7482_/A sky130_fd_sc_hd__o22a_1
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9218_ _9823_/Q _7649_/Y _9528_/Q vssd1 vssd1 vccd1 vccd1 _9218_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9149_ _6190_/Y input17/X _9155_/S vssd1 vssd1 vccd1 vccd1 _9149_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6850_ _6847_/A _6847_/B _6847_/X vssd1 vssd1 vccd1 vccd1 _6851_/B sky130_fd_sc_hd__a21bo_1
X_5801_ _5801_/A vssd1 vssd1 vccd1 vccd1 _7086_/A sky130_fd_sc_hd__inv_2
XFILLER_50_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6781_ _6781_/A _6787_/A vssd1 vssd1 vccd1 vccd1 _6781_/Y sky130_fd_sc_hd__nor2_1
X_8520_ _8483_/X _8519_/X _8483_/X _8519_/X vssd1 vssd1 vccd1 vccd1 _8521_/A sky130_fd_sc_hd__a2bb2o_2
X_5732_ _9674_/Q _9657_/Q vssd1 vssd1 vccd1 vccd1 _5732_/Y sky130_fd_sc_hd__nor2_1
XFILLER_200_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8451_ _8475_/C _8436_/X _8426_/A vssd1 vssd1 vccd1 vccd1 _8455_/A sky130_fd_sc_hd__a21oi_2
XFILLER_148_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5663_ _9688_/Q _5658_/X _9672_/Q _5662_/X _5660_/X vssd1 vssd1 vccd1 vccd1 _9688_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_209_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5594_ _5594_/A vssd1 vssd1 vccd1 vccd1 _5594_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8382_ _9696_/Q _6596_/Y _9696_/Q _6596_/Y vssd1 vssd1 vccd1 vccd1 _8382_/X sky130_fd_sc_hd__a2bb2o_1
X_7402_ _7384_/A _7384_/B _7384_/C _7407_/B vssd1 vssd1 vccd1 vccd1 _7403_/A sky130_fd_sc_hd__o22a_1
XFILLER_190_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7333_ _7325_/X _7326_/X _7325_/X _7326_/X vssd1 vssd1 vccd1 vccd1 _7351_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_116_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9003_ _9780_/Q _9897_/Q _9480_/S vssd1 vssd1 vccd1 vccd1 _9003_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7264_ _7290_/A _9469_/X vssd1 vssd1 vccd1 vccd1 _7264_/X sky130_fd_sc_hd__or2_1
X_7195_ _7195_/A vssd1 vssd1 vccd1 vccd1 _7201_/A sky130_fd_sc_hd__clkbuf_2
X_6215_ _9578_/Q vssd1 vssd1 vccd1 vccd1 _8010_/A sky130_fd_sc_hd__inv_2
XFILLER_112_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6146_ _6146_/A vssd1 vssd1 vccd1 vccd1 _6165_/A sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_14 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6077_ _7986_/A _9645_/Q _6066_/A _6068_/Y vssd1 vssd1 vccd1 vccd1 _6077_/X sky130_fd_sc_hd__a22o_1
X_5028_ _5028_/A vssd1 vssd1 vccd1 vccd1 _5028_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_9905_ _9917_/CLK _9905_/D vssd1 vssd1 vccd1 vccd1 _9905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9836_ _9836_/CLK _9836_/D vssd1 vssd1 vccd1 vccd1 _9836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6979_ _6682_/X _6685_/X _6681_/X vssd1 vssd1 vccd1 vccd1 _6979_/X sky130_fd_sc_hd__o21a_1
X_9767_ _9916_/CLK _9767_/D vssd1 vssd1 vccd1 vccd1 _9767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8718_ _8713_/X _8717_/Y _8713_/X _8717_/Y vssd1 vssd1 vccd1 vccd1 _8718_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_139_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9698_ _9699_/CLK _9698_/D vssd1 vssd1 vccd1 vccd1 _9698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8649_ _8650_/B vssd1 vssd1 vccd1 vccd1 _8649_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6000_ _5998_/X _5999_/Y _5998_/X _5999_/Y vssd1 vssd1 vccd1 vccd1 _6000_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_39_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7951_ _8630_/A vssd1 vssd1 vccd1 vccd1 _8776_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7882_ _7882_/A _7882_/B vssd1 vssd1 vccd1 vccd1 _7887_/B sky130_fd_sc_hd__or2_1
XFILLER_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6902_ _6902_/A _6902_/B vssd1 vssd1 vccd1 vccd1 _6903_/B sky130_fd_sc_hd__or2_1
XFILLER_211_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9621_ _9715_/CLK _9621_/D vssd1 vssd1 vccd1 vccd1 _9621_/Q sky130_fd_sc_hd__dfxtp_1
X_6833_ _6833_/A _6833_/B vssd1 vssd1 vccd1 vccd1 _6834_/B sky130_fd_sc_hd__or2_2
XFILLER_35_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9552_ _9923_/CLK _9552_/D vssd1 vssd1 vccd1 vccd1 _9552_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6764_ _6764_/A _6764_/B vssd1 vssd1 vccd1 vccd1 _6765_/A sky130_fd_sc_hd__or2_4
XFILLER_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8503_ _8534_/A _9378_/X _8472_/A _8625_/B vssd1 vssd1 vccd1 vccd1 _8503_/X sky130_fd_sc_hd__o22a_1
X_5715_ _9681_/Q _9664_/Q vssd1 vssd1 vccd1 vccd1 _5715_/Y sky130_fd_sc_hd__nor2_1
X_9483_ _9482_/X _8935_/A _9505_/S vssd1 vssd1 vccd1 vccd1 _9483_/X sky130_fd_sc_hd__mux2_1
X_6695_ _6867_/D vssd1 vssd1 vccd1 vccd1 _6883_/A sky130_fd_sc_hd__clkbuf_2
X_8434_ _8471_/A _8469_/B vssd1 vssd1 vccd1 vccd1 _8472_/C sky130_fd_sc_hd__nor2_4
X_5646_ _9678_/Q vssd1 vssd1 vccd1 vccd1 _6577_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8365_ _8357_/B _8356_/X _8360_/X vssd1 vssd1 vccd1 vccd1 _8365_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_191_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5577_ _8967_/B vssd1 vssd1 vccd1 vccd1 _5577_/X sky130_fd_sc_hd__clkbuf_2
X_8296_ _7897_/A _8202_/X _7902_/A _8201_/Y _8295_/X vssd1 vssd1 vccd1 vccd1 _8296_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_116_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7316_ _7314_/X _7315_/X _7314_/X _7315_/X vssd1 vssd1 vccd1 vccd1 _7323_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7247_ _7247_/A _7247_/B vssd1 vssd1 vccd1 vccd1 _7259_/A sky130_fd_sc_hd__or2_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7178_ _7178_/A _7178_/B vssd1 vssd1 vccd1 vccd1 _7190_/A sky130_fd_sc_hd__or2_1
XFILLER_105_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6129_ _9564_/Q _6146_/A _9563_/Q _6123_/X vssd1 vssd1 vccd1 vccd1 _6130_/B sky130_fd_sc_hd__a22o_1
XFILLER_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9819_ _9819_/CLK _9819_/D vssd1 vssd1 vccd1 vccd1 _9819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5500_ _9416_/X _5499_/X _9416_/X _5499_/X vssd1 vssd1 vccd1 vccd1 _5600_/A sky130_fd_sc_hd__a2bb2oi_1
XFILLER_13_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6480_ _6480_/A _6480_/B _6480_/C vssd1 vssd1 vccd1 vccd1 _6480_/X sky130_fd_sc_hd__or3_1
XFILLER_118_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5431_ _5431_/A _5431_/B vssd1 vssd1 vccd1 vccd1 _5431_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8150_ _7698_/X _8114_/X _8149_/Y vssd1 vssd1 vccd1 vccd1 _8150_/X sky130_fd_sc_hd__o21ba_1
X_5362_ _9726_/Q _5362_/B vssd1 vssd1 vccd1 vccd1 _5362_/Y sky130_fd_sc_hd__nor2_1
X_8081_ _9553_/Q _8081_/B vssd1 vssd1 vccd1 vccd1 _8082_/B sky130_fd_sc_hd__or2_1
XFILLER_160_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7101_ _7407_/B vssd1 vssd1 vccd1 vccd1 _7101_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_141_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5293_ _5293_/A vssd1 vssd1 vccd1 vccd1 _9738_/D sky130_fd_sc_hd__inv_2
X_7032_ _7022_/X _7023_/X _7024_/X _7031_/X vssd1 vssd1 vccd1 vccd1 _7032_/X sky130_fd_sc_hd__o22a_1
XFILLER_82_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8983_ _8982_/X _7490_/A _9506_/S vssd1 vssd1 vccd1 vccd1 _8983_/X sky130_fd_sc_hd__mux2_1
X_7934_ _8821_/A vssd1 vssd1 vccd1 vccd1 _8938_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7865_ _7865_/A _7865_/B vssd1 vssd1 vccd1 vccd1 _7869_/B sky130_fd_sc_hd__or2_1
XPHY_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7796_ _8123_/A _7659_/B _7795_/Y vssd1 vssd1 vccd1 vccd1 _7796_/X sky130_fd_sc_hd__a21o_1
XPHY_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6816_ _6586_/A _9427_/X _6796_/C _6796_/D vssd1 vssd1 vccd1 vccd1 _6817_/A sky130_fd_sc_hd__o22a_1
XPHY_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9604_ _9895_/CLK _9604_/D vssd1 vssd1 vccd1 vccd1 _9604_/Q sky130_fd_sc_hd__dfxtp_1
X_9535_ _9796_/CLK _9535_/D vssd1 vssd1 vccd1 vccd1 _9535_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6747_ _6764_/A _6760_/B _6814_/A _6764_/B vssd1 vssd1 vccd1 vccd1 _6749_/A sky130_fd_sc_hd__o22a_1
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9466_ _6596_/Y _6597_/Y _9683_/Q vssd1 vssd1 vccd1 vccd1 _9466_/X sky130_fd_sc_hd__mux2_1
X_6678_ _6678_/A vssd1 vssd1 vccd1 vccd1 _6978_/A sky130_fd_sc_hd__buf_2
X_8417_ _8469_/B vssd1 vssd1 vccd1 vccd1 _8543_/B sky130_fd_sc_hd__buf_2
X_5629_ _5704_/A _5626_/Y _5627_/X _7636_/A _5607_/X vssd1 vssd1 vccd1 vccd1 _5630_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_136_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9397_ _9795_/Q _9912_/Q _9480_/S vssd1 vssd1 vccd1 vccd1 _9397_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8348_ _8340_/B _8339_/X _8343_/X vssd1 vssd1 vccd1 vccd1 _8348_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8279_ _7715_/X _8228_/Y _8278_/X vssd1 vssd1 vccd1 vccd1 _8279_/X sky130_fd_sc_hd__a21o_1
XFILLER_116_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5980_ _7928_/A _9636_/Q _9849_/Q _5979_/Y vssd1 vssd1 vccd1 vccd1 _5981_/A sky130_fd_sc_hd__o22a_1
XFILLER_37_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4931_ _5815_/A _5815_/B _4931_/C _5881_/A vssd1 vssd1 vccd1 vccd1 _5967_/A sky130_fd_sc_hd__or4_4
X_7650_ _7650_/A _7652_/B vssd1 vssd1 vccd1 vccd1 _7650_/Y sky130_fd_sc_hd__nor2_1
X_4862_ _9896_/Q vssd1 vssd1 vccd1 vccd1 _5222_/A sky130_fd_sc_hd__inv_2
XFILLER_205_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6601_ _6867_/A vssd1 vssd1 vccd1 vccd1 _6890_/B sky130_fd_sc_hd__buf_1
XFILLER_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9320_ _9776_/Q _9319_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9320_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4793_ _9919_/Q vssd1 vssd1 vccd1 vccd1 _4794_/A sky130_fd_sc_hd__clkbuf_2
X_7581_ _7581_/A vssd1 vssd1 vccd1 vccd1 _7601_/A sky130_fd_sc_hd__inv_2
XFILLER_158_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6532_ _6535_/A _6532_/B vssd1 vssd1 vccd1 vccd1 _6532_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9251_ _7806_/X _9755_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9251_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6463_ _6463_/A _6463_/B _6463_/C _6462_/X vssd1 vssd1 vccd1 vccd1 _6463_/X sky130_fd_sc_hd__or4b_4
XFILLER_9_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8202_ _8200_/A _8200_/B _8200_/Y vssd1 vssd1 vccd1 vccd1 _8202_/X sky130_fd_sc_hd__a21o_1
XFILLER_133_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9182_ _6521_/Y _9787_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9536_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5414_ _9356_/X vssd1 vssd1 vccd1 vccd1 _5415_/B sky130_fd_sc_hd__inv_2
X_6394_ _9776_/Q _8199_/A vssd1 vssd1 vccd1 vccd1 _6402_/A sky130_fd_sc_hd__or2_1
X_8133_ _7749_/A _8128_/X _9899_/Q _8131_/Y _8132_/X vssd1 vssd1 vccd1 vccd1 _8133_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_99_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5345_ _5337_/A _5341_/Y _5344_/Y _5340_/X vssd1 vssd1 vccd1 vccd1 _9730_/D sky130_fd_sc_hd__a2bb2o_1
X_8064_ _9536_/Q _8064_/B vssd1 vssd1 vccd1 vccd1 _8065_/B sky130_fd_sc_hd__or2_1
XFILLER_99_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5276_ _5268_/B _5271_/X _5273_/Y _5275_/X _5247_/A vssd1 vssd1 vccd1 vccd1 _5277_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_101_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7015_ _7013_/X _7014_/X _7013_/X _7014_/X vssd1 vssd1 vccd1 vccd1 _7015_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8966_ _8931_/X _8965_/Y _8931_/X _8965_/Y vssd1 vssd1 vccd1 vccd1 _8966_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_102_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7917_ _9507_/X _8378_/A vssd1 vssd1 vccd1 vccd1 _7917_/X sky130_fd_sc_hd__and2_1
XFILLER_70_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8897_ _8897_/A vssd1 vssd1 vccd1 vccd1 _8897_/Y sky130_fd_sc_hd__inv_2
XPHY_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7848_ _7848_/A _7848_/B vssd1 vssd1 vccd1 vccd1 _7852_/B sky130_fd_sc_hd__or2_1
XPHY_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7779_ _7779_/A _7783_/B vssd1 vssd1 vccd1 vccd1 _7780_/A sky130_fd_sc_hd__or2_1
XPHY_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9518_ _9907_/CLK _9518_/D vssd1 vssd1 vccd1 vccd1 _9518_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9449_ _6334_/Y _7761_/X _9480_/S vssd1 vssd1 vccd1 vccd1 _9449_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 io_wb_adr_i[8] vssd1 vssd1 vccd1 vccd1 _4855_/A sky130_fd_sc_hd__buf_1
XFILLER_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput35 io_wb_dat_i[27] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_4
Xinput24 io_wb_dat_i[17] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_4
XPHY_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput46 io_wb_dat_i[8] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_6
XFILLER_115_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5130_ _5138_/A vssd1 vssd1 vccd1 vccd1 _5130_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5061_ _5136_/A vssd1 vssd1 vccd1 vccd1 _5061_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8820_ _8944_/C _8942_/B vssd1 vssd1 vccd1 vccd1 _8820_/X sky130_fd_sc_hd__or2_2
XFILLER_80_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8751_ _8942_/A _8751_/B _8823_/C vssd1 vssd1 vccd1 vccd1 _8751_/X sky130_fd_sc_hd__or3_4
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5963_ _9143_/X _5958_/X _9566_/Q _5959_/X vssd1 vssd1 vccd1 vccd1 _9566_/D sky130_fd_sc_hd__a22o_1
XFILLER_178_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7702_ _9917_/Q vssd1 vssd1 vccd1 vccd1 _7861_/A sky130_fd_sc_hd__inv_2
X_4914_ _5631_/A vssd1 vssd1 vccd1 vccd1 _4914_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8682_ _8680_/X _8681_/X _8680_/X _8681_/X vssd1 vssd1 vccd1 vccd1 _8682_/X sky130_fd_sc_hd__a2bb2o_1
X_5894_ _9613_/Q _5884_/A _4860_/A _5885_/A _5891_/X vssd1 vssd1 vccd1 vccd1 _9613_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4845_ _4923_/A vssd1 vssd1 vccd1 vccd1 _4845_/X sky130_fd_sc_hd__clkbuf_4
X_7633_ _7487_/A _7101_/X _7577_/X _7591_/A vssd1 vssd1 vccd1 vccd1 _7633_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_119_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4776_ _4776_/A vssd1 vssd1 vccd1 vccd1 _5405_/A sky130_fd_sc_hd__clkbuf_2
X_7564_ _7603_/A vssd1 vssd1 vccd1 vccd1 _7564_/Y sky130_fd_sc_hd__inv_2
X_6515_ _9808_/Q _6547_/B _9809_/Q _6548_/B _6514_/X vssd1 vssd1 vccd1 vccd1 _6515_/Y
+ sky130_fd_sc_hd__o221ai_1
X_9303_ _7876_/Y _9772_/Q _9327_/S vssd1 vssd1 vccd1 vccd1 _9303_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7495_ _7493_/Y _7494_/X _7493_/Y _7494_/X vssd1 vssd1 vccd1 vccd1 _7495_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_173_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9234_ _9233_/X _4860_/A _9334_/S vssd1 vssd1 vccd1 vccd1 _9234_/X sky130_fd_sc_hd__mux2_1
X_6446_ _9788_/Q _6522_/B _6338_/Y _6447_/A vssd1 vssd1 vccd1 vccd1 _6446_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_106_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9165_ _6278_/X input34/X _9170_/S vssd1 vssd1 vccd1 vccd1 _9165_/X sky130_fd_sc_hd__mux2_1
X_6377_ _9759_/Q _6377_/B vssd1 vssd1 vccd1 vccd1 _8231_/A sky130_fd_sc_hd__or2_2
XFILLER_161_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8116_ _9540_/Q _8068_/B _8069_/B vssd1 vssd1 vccd1 vccd1 _8116_/X sky130_fd_sc_hd__a21bo_1
XFILLER_88_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9096_ _5982_/X _5983_/X _9896_/Q vssd1 vssd1 vccd1 vccd1 _9096_/X sky130_fd_sc_hd__mux2_1
X_5328_ _5328_/A _5384_/A vssd1 vssd1 vccd1 vccd1 _5380_/A sky130_fd_sc_hd__or2_1
X_8047_ _9448_/X _8047_/B vssd1 vssd1 vccd1 vccd1 _8047_/X sky130_fd_sc_hd__and2_1
XFILLER_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5259_ _5259_/A vssd1 vssd1 vccd1 vccd1 _5260_/B sky130_fd_sc_hd__inv_2
XFILLER_68_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8949_ _8937_/X _8948_/X _8937_/X _8948_/X vssd1 vssd1 vccd1 vccd1 _8949_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_71_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6300_ _8044_/A _6193_/A _6295_/X _6297_/X vssd1 vssd1 vccd1 vccd1 _6300_/X sky130_fd_sc_hd__o22a_1
XFILLER_116_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clock/X
+ sky130_fd_sc_hd__clkbuf_1
X_7280_ _7266_/Y _7267_/X _7278_/X _7279_/X vssd1 vssd1 vccd1 vccd1 _7280_/X sky130_fd_sc_hd__o22a_1
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6231_ _9581_/Q _6169_/A _8017_/A _6139_/A vssd1 vssd1 vccd1 vccd1 _6244_/A sky130_fd_sc_hd__a22o_1
XFILLER_131_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6162_ _6159_/X _6161_/Y _6159_/X _6161_/Y vssd1 vssd1 vccd1 vccd1 _6162_/X sky130_fd_sc_hd__o2bb2a_1
X_5113_ _9829_/Q vssd1 vssd1 vccd1 vccd1 _5113_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6093_ _9648_/Q vssd1 vssd1 vccd1 vccd1 _6094_/B sky130_fd_sc_hd__inv_2
X_5044_ _5070_/A vssd1 vssd1 vccd1 vccd1 _5069_/A sky130_fd_sc_hd__clkbuf_2
X_9921_ _9923_/CLK _9921_/D vssd1 vssd1 vccd1 vccd1 _9921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9852_ _9879_/CLK _9852_/D vssd1 vssd1 vccd1 vccd1 _9852_/Q sky130_fd_sc_hd__dfxtp_2
X_8803_ _8803_/A vssd1 vssd1 vccd1 vccd1 _8803_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9783_ _9819_/CLK _9783_/D vssd1 vssd1 vccd1 vccd1 _9783_/Q sky130_fd_sc_hd__dfxtp_1
X_6995_ _6995_/A _6995_/B vssd1 vssd1 vccd1 vccd1 _6995_/X sky130_fd_sc_hd__or2_1
XFILLER_25_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8734_ _8755_/A _9395_/X vssd1 vssd1 vccd1 vccd1 _8734_/X sky130_fd_sc_hd__or2_2
XFILLER_80_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5946_ _9155_/X _5944_/X _9579_/Q _5945_/X vssd1 vssd1 vccd1 vccd1 _9579_/D sky130_fd_sc_hd__a22o_1
XFILLER_40_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8665_ _8709_/B vssd1 vssd1 vccd1 vccd1 _8665_/Y sky130_fd_sc_hd__inv_2
X_5877_ _9620_/Q vssd1 vssd1 vccd1 vccd1 _7273_/A sky130_fd_sc_hd__clkbuf_2
X_4828_ _9905_/Q vssd1 vssd1 vccd1 vccd1 _7810_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7616_ _7076_/A _7076_/B _7077_/B vssd1 vssd1 vccd1 vccd1 _7616_/X sky130_fd_sc_hd__a21bo_1
X_8596_ _8596_/A _8596_/B vssd1 vssd1 vccd1 vccd1 _8596_/Y sky130_fd_sc_hd__nor2_8
XFILLER_21_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4759_ _4743_/X _4753_/Y _4753_/A _4754_/X _5916_/A vssd1 vssd1 vccd1 vccd1 _9929_/D
+ sky130_fd_sc_hd__o221a_1
X_7547_ _7457_/X _7470_/Y _7471_/X _7473_/A vssd1 vssd1 vccd1 vccd1 _7548_/B sky130_fd_sc_hd__a31o_1
XFILLER_175_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7478_ _7437_/X _7476_/X _7537_/B vssd1 vssd1 vccd1 vccd1 _7478_/X sky130_fd_sc_hd__o21a_1
XFILLER_161_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9217_ _9822_/Q _7648_/Y _9528_/Q vssd1 vssd1 vccd1 vccd1 _9217_/X sky130_fd_sc_hd__mux2_1
X_6429_ _9763_/Q vssd1 vssd1 vccd1 vccd1 _6429_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9148_ _6184_/X input47/X _9148_/S vssd1 vssd1 vccd1 vccd1 _9148_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9079_ _9078_/X input20/X _9282_/S vssd1 vssd1 vccd1 vccd1 _9079_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5800_ _5739_/X _5746_/X _5739_/X _5746_/X vssd1 vssd1 vccd1 vccd1 _5801_/A sky130_fd_sc_hd__a2bb2o_1
X_6780_ _6765_/A _6775_/Y _6772_/X _6776_/X vssd1 vssd1 vccd1 vccd1 _6787_/A sky130_fd_sc_hd__o22ai_4
XFILLER_35_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5731_ _9675_/Q _9658_/Q vssd1 vssd1 vccd1 vccd1 _5731_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8450_ _8499_/A _8450_/B vssd1 vssd1 vccd1 vccd1 _8457_/A sky130_fd_sc_hd__or2_1
X_5662_ _5662_/A vssd1 vssd1 vccd1 vccd1 _5662_/X sky130_fd_sc_hd__clkbuf_2
X_8381_ _8381_/A _8381_/B vssd1 vssd1 vccd1 vccd1 _8381_/Y sky130_fd_sc_hd__nor2_1
X_5593_ _9707_/Q _4922_/X _5570_/X _5592_/Y _5187_/X vssd1 vssd1 vccd1 vccd1 _9707_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7401_ _7397_/X _7400_/X _7397_/X _7400_/X vssd1 vssd1 vccd1 vccd1 _7401_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_209_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7332_ _7327_/X _7331_/X _7327_/X _7331_/X vssd1 vssd1 vccd1 vccd1 _7332_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_143_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7263_ _7241_/X _7262_/X _7241_/X _7262_/X vssd1 vssd1 vccd1 vccd1 _7263_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_171_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9002_ _9001_/X _6352_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _9002_/X sky130_fd_sc_hd__mux2_1
X_6214_ _6221_/C _6213_/X _6221_/C _6213_/X vssd1 vssd1 vccd1 vccd1 _6214_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_171_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7194_ _7172_/X _7193_/X _7172_/X _7193_/X vssd1 vssd1 vccd1 vccd1 _7194_/X sky130_fd_sc_hd__a2bb2o_1
X_6145_ _6150_/B _6144_/Y _6150_/B _6144_/Y vssd1 vssd1 vccd1 vccd1 _6145_/X sky130_fd_sc_hd__a2bb2o_1
XINSDIODE2_15 input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6076_ _6076_/A vssd1 vssd1 vccd1 vccd1 _6076_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5027_ _9819_/Q _5019_/X _5026_/X _5020_/X _5024_/X vssd1 vssd1 vccd1 vccd1 _9819_/D
+ sky130_fd_sc_hd__o221a_1
X_9904_ _9917_/CLK _9904_/D vssd1 vssd1 vccd1 vccd1 _9904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9835_ _9836_/CLK _9835_/D vssd1 vssd1 vccd1 vccd1 _9835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_32_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _9761_/CLK sky130_fd_sc_hd__clkbuf_16
X_9766_ _9916_/CLK _9766_/D vssd1 vssd1 vccd1 vccd1 _9766_/Q sky130_fd_sc_hd__dfxtp_1
X_8717_ _8717_/A vssd1 vssd1 vccd1 vccd1 _8717_/Y sky130_fd_sc_hd__inv_2
X_6978_ _6978_/A _9465_/X _6978_/C _9466_/X vssd1 vssd1 vccd1 vccd1 _6978_/X sky130_fd_sc_hd__or4_4
XFILLER_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5929_ _9166_/X _5921_/X _9590_/Q _5924_/X vssd1 vssd1 vccd1 vccd1 _9590_/D sky130_fd_sc_hd__a22o_1
XFILLER_139_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9697_ _9697_/CLK _9697_/D vssd1 vssd1 vccd1 vccd1 _9697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8648_ _8405_/Y _8647_/X _8405_/Y _8647_/X vssd1 vssd1 vccd1 vccd1 _8650_/B sky130_fd_sc_hd__a2bb2o_1
X_8579_ _8561_/X _8578_/X _8561_/X _8578_/X vssd1 vssd1 vccd1 vccd1 _8593_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_119_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7950_ _9632_/Q vssd1 vssd1 vccd1 vccd1 _8630_/A sky130_fd_sc_hd__inv_2
XFILLER_94_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7881_ _7882_/A vssd1 vssd1 vccd1 vccd1 _7881_/X sky130_fd_sc_hd__buf_2
XFILLER_94_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6901_ _6877_/C _6874_/B _6874_/Y vssd1 vssd1 vccd1 vccd1 _6902_/B sky130_fd_sc_hd__o21ai_1
XFILLER_211_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6832_ _6807_/C _6803_/X _6807_/C _6803_/X vssd1 vssd1 vccd1 vccd1 _6833_/B sky130_fd_sc_hd__o2bb2ai_1
X_9620_ _9715_/CLK _9620_/D vssd1 vssd1 vccd1 vccd1 _9620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9551_ _9923_/CLK _9551_/D vssd1 vssd1 vccd1 vccd1 _9551_/Q sky130_fd_sc_hd__dfxtp_1
X_6763_ _6749_/X _6750_/X _6761_/X _6762_/X vssd1 vssd1 vccd1 vccd1 _6763_/X sky130_fd_sc_hd__o22a_1
XFILLER_195_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8502_ _9377_/X vssd1 vssd1 vccd1 vccd1 _8625_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_188_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5714_ _6982_/A _9665_/Q _6598_/A _5713_/Y vssd1 vssd1 vccd1 vccd1 _5714_/X sky130_fd_sc_hd__a22o_1
X_9482_ _7928_/X _5979_/Y _9504_/S vssd1 vssd1 vccd1 vccd1 _9482_/X sky130_fd_sc_hd__mux2_1
X_6694_ _9618_/Q vssd1 vssd1 vccd1 vccd1 _6867_/D sky130_fd_sc_hd__inv_2
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8433_ _8431_/Y _8430_/X _8446_/A vssd1 vssd1 vccd1 vccd1 _8433_/Y sky130_fd_sc_hd__o21ai_1
X_5645_ _5689_/A vssd1 vssd1 vccd1 vccd1 _5645_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8364_ _8347_/X _8351_/X _8375_/C vssd1 vssd1 vccd1 vccd1 _8364_/X sky130_fd_sc_hd__o21ba_1
X_5576_ _5644_/A vssd1 vssd1 vccd1 vccd1 _8967_/B sky130_fd_sc_hd__buf_2
X_8295_ _7897_/A _8202_/X _7892_/A _8206_/X _8294_/X vssd1 vssd1 vccd1 vccd1 _8295_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7315_ _7324_/A _9474_/X vssd1 vssd1 vccd1 vccd1 _7315_/X sky130_fd_sc_hd__or2_1
XFILLER_171_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7246_ _7233_/X _7234_/X _7233_/X _7234_/X vssd1 vssd1 vccd1 vccd1 _7246_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7177_ _7164_/X _7165_/X _7164_/X _7165_/X vssd1 vssd1 vccd1 vccd1 _7177_/X sky130_fd_sc_hd__a2bb2o_2
X_6128_ _6125_/Y _6148_/A _9565_/Q _6146_/A vssd1 vssd1 vccd1 vccd1 _6130_/A sky130_fd_sc_hd__o22a_1
XFILLER_58_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6059_ _6059_/A vssd1 vssd1 vccd1 vccd1 _6059_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9818_ _9929_/CLK _9818_/D vssd1 vssd1 vccd1 vccd1 _9818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9749_ _9750_/CLK _9749_/D vssd1 vssd1 vccd1 vccd1 _9749_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_41_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5430_ _9341_/X vssd1 vssd1 vccd1 vccd1 _5431_/B sky130_fd_sc_hd__inv_2
XFILLER_173_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5361_ _5361_/A vssd1 vssd1 vccd1 vccd1 _5362_/B sky130_fd_sc_hd__inv_2
X_8080_ _9552_/Q _8080_/B vssd1 vssd1 vccd1 vccd1 _8081_/B sky130_fd_sc_hd__or2_4
XFILLER_113_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5292_ _5287_/B _5271_/X _5291_/Y _5275_/X _5243_/A vssd1 vssd1 vccd1 vccd1 _5293_/A
+ sky130_fd_sc_hd__o32a_1
X_7100_ _7389_/B vssd1 vssd1 vccd1 vccd1 _7407_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_113_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7031_ _7025_/X _7027_/X _7028_/X _7030_/X vssd1 vssd1 vccd1 vccd1 _7031_/X sky130_fd_sc_hd__o22a_1
XFILLER_141_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8982_ _8981_/X _8955_/A _9505_/S vssd1 vssd1 vccd1 vccd1 _8982_/X sky130_fd_sc_hd__mux2_1
X_7933_ _8534_/A vssd1 vssd1 vccd1 vccd1 _8821_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7864_ _4798_/X _7675_/B _7863_/Y vssd1 vssd1 vccd1 vccd1 _7864_/X sky130_fd_sc_hd__a21o_1
XPHY_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7795_ _7795_/A vssd1 vssd1 vccd1 vccd1 _7795_/Y sky130_fd_sc_hd__inv_2
XPHY_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9603_ _9895_/CLK _9603_/D vssd1 vssd1 vccd1 vccd1 _9603_/Q sky130_fd_sc_hd__dfxtp_1
X_6815_ _6810_/X _6814_/X _6810_/X _6814_/X vssd1 vssd1 vccd1 vccd1 _6815_/X sky130_fd_sc_hd__a2bb2o_1
X_9534_ _9796_/CLK _9534_/D vssd1 vssd1 vccd1 vccd1 _9534_/Q sky130_fd_sc_hd__dfxtp_1
X_6746_ _6724_/X _6745_/X _6724_/X _6745_/X vssd1 vssd1 vccd1 vccd1 _6746_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9465_ _6591_/Y _6595_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9465_/X sky130_fd_sc_hd__mux2_2
X_6677_ _9466_/X vssd1 vssd1 vccd1 vccd1 _6981_/B sky130_fd_sc_hd__buf_1
X_8416_ _8416_/A vssd1 vssd1 vccd1 vccd1 _8469_/B sky130_fd_sc_hd__clkbuf_2
X_5628_ _9700_/Q vssd1 vssd1 vccd1 vccd1 _7636_/A sky130_fd_sc_hd__inv_2
X_9396_ _8748_/Y _8747_/B _9477_/S vssd1 vssd1 vccd1 vccd1 _9396_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8347_ _8316_/X _8332_/Y _8375_/D vssd1 vssd1 vccd1 vccd1 _8347_/X sky130_fd_sc_hd__o21ba_1
X_5559_ _5579_/A _5559_/B vssd1 vssd1 vccd1 vccd1 _9714_/D sky130_fd_sc_hd__nor2_1
XFILLER_105_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8278_ _7713_/X _8230_/X _7840_/A _8228_/Y _8277_/X vssd1 vssd1 vccd1 vccd1 _8278_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_132_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7229_ _7385_/A _7359_/A vssd1 vssd1 vccd1 vccd1 _7230_/C sky130_fd_sc_hd__or2_1
XFILLER_116_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4930_ _5917_/A _5862_/A vssd1 vssd1 vccd1 vccd1 _5881_/A sky130_fd_sc_hd__or2_1
X_4861_ _4853_/X _8999_/S _4860_/X _4859_/A _4845_/X vssd1 vssd1 vccd1 vccd1 _9896_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_45_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6600_ _9617_/Q vssd1 vssd1 vccd1 vccd1 _6867_/A sky130_fd_sc_hd__inv_2
XFILLER_165_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4792_ _9087_/X _4782_/X _4790_/X _4784_/X _4791_/X vssd1 vssd1 vccd1 vccd1 _9920_/D
+ sky130_fd_sc_hd__o221a_1
X_7580_ _7580_/A vssd1 vssd1 vccd1 vccd1 _7602_/A sky130_fd_sc_hd__inv_2
X_6531_ _6535_/A _6531_/B vssd1 vssd1 vccd1 vccd1 _6531_/Y sky130_fd_sc_hd__nor2_1
X_9250_ _9249_/X _5029_/A _9306_/S vssd1 vssd1 vccd1 vccd1 _9250_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6462_ _6451_/Y _6462_/B _6462_/C _6462_/D vssd1 vssd1 vccd1 vccd1 _6462_/X sky130_fd_sc_hd__and4b_1
X_6393_ _9775_/Q _6393_/B vssd1 vssd1 vccd1 vccd1 _8199_/A sky130_fd_sc_hd__or2_2
X_8201_ _6343_/Y _8200_/Y _8197_/Y vssd1 vssd1 vccd1 vccd1 _8201_/Y sky130_fd_sc_hd__o21bai_1
X_9181_ _6520_/Y _9786_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9535_/D sky130_fd_sc_hd__mux2_1
X_5413_ _9360_/X vssd1 vssd1 vccd1 vccd1 _5415_/A sky130_fd_sc_hd__inv_2
X_8132_ _8057_/A _8057_/B _9898_/Q _8128_/X _8057_/Y vssd1 vssd1 vccd1 vccd1 _8132_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5344_ _5344_/A vssd1 vssd1 vccd1 vccd1 _5344_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8063_ _9535_/Q _8063_/B vssd1 vssd1 vccd1 vccd1 _8064_/B sky130_fd_sc_hd__or2_1
XFILLER_87_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5275_ _5275_/A vssd1 vssd1 vccd1 vccd1 _5275_/X sky130_fd_sc_hd__clkbuf_2
X_7014_ _7003_/A _7003_/B _7003_/X vssd1 vssd1 vccd1 vccd1 _7014_/X sky130_fd_sc_hd__a21bo_1
XFILLER_68_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8965_ _8949_/X _8964_/X _8949_/X _8964_/X vssd1 vssd1 vccd1 vccd1 _8965_/Y sky130_fd_sc_hd__a2bb2oi_4
XFILLER_55_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8896_ _8811_/A _8812_/A _8857_/Y _8854_/Y _8895_/X vssd1 vssd1 vccd1 vccd1 _8897_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_102_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7916_ _7991_/A vssd1 vssd1 vccd1 vccd1 _8378_/A sky130_fd_sc_hd__inv_2
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7847_ _9914_/Q _7671_/B _7846_/Y vssd1 vssd1 vccd1 vccd1 _7847_/X sky130_fd_sc_hd__a21o_1
XPHY_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7778_ _8322_/A _7778_/B vssd1 vssd1 vccd1 vccd1 _7783_/B sky130_fd_sc_hd__nor2_2
XPHY_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9517_ _9519_/CLK _9517_/D vssd1 vssd1 vccd1 vccd1 _9518_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_149_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6729_ _6716_/X _6717_/X _6716_/X _6717_/X vssd1 vssd1 vccd1 vccd1 _6729_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9448_ _9447_/X _9779_/Q _9481_/S vssd1 vssd1 vccd1 vccd1 _9448_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9379_ _8419_/Y _8415_/X _9477_/S vssd1 vssd1 vccd1 vccd1 _9379_/X sky130_fd_sc_hd__mux2_4
XFILLER_152_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput36 io_wb_dat_i[28] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_4
Xinput25 io_wb_dat_i[18] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_4
XPHY_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 io_wb_adr_i[9] vssd1 vssd1 vccd1 vccd1 _4856_/C sky130_fd_sc_hd__buf_1
XFILLER_155_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput47 io_wb_dat_i[9] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__buf_6
XFILLER_182_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5060_ _5069_/A _5060_/B vssd1 vssd1 vccd1 vccd1 _9809_/D sky130_fd_sc_hd__nor2_1
XFILLER_69_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8750_ _8938_/A _8751_/B _8865_/A _8875_/D vssd1 vssd1 vccd1 vccd1 _8752_/A sky130_fd_sc_hd__o22a_1
XFILLER_25_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5962_ _9144_/X _5958_/X _9567_/Q _5959_/X vssd1 vssd1 vccd1 vccd1 _9567_/D sky130_fd_sc_hd__a22o_1
XFILLER_206_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7701_ _7696_/X _5198_/X _7698_/X _9761_/Q _7700_/X vssd1 vssd1 vccd1 vccd1 _7705_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_92_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4913_ _9872_/Q _4905_/X _9724_/Q _4912_/X _4906_/X vssd1 vssd1 vccd1 vccd1 _9872_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8681_ _8624_/X _8635_/X _8637_/A _8638_/A vssd1 vssd1 vccd1 vccd1 _8681_/X sky130_fd_sc_hd__o22a_1
X_5893_ _9614_/Q _5884_/A _5035_/A _5885_/A _5891_/X vssd1 vssd1 vccd1 vccd1 _9614_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_166_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7632_ _6573_/X _6982_/D _7055_/X _7068_/A vssd1 vssd1 vccd1 vccd1 _7632_/Y sky130_fd_sc_hd__o31ai_1
X_4844_ _5405_/A vssd1 vssd1 vccd1 vccd1 _4923_/A sky130_fd_sc_hd__buf_2
XFILLER_21_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4775_ _7682_/A vssd1 vssd1 vccd1 vccd1 _4775_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7563_ _7552_/Y _7562_/Y _7552_/Y _7562_/Y vssd1 vssd1 vccd1 vccd1 _7603_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_193_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6514_ _9808_/Q _6547_/B _9807_/Q _6546_/B _6513_/X vssd1 vssd1 vccd1 vccd1 _6514_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_165_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9302_ _9301_/X input30/X _9306_/S vssd1 vssd1 vccd1 vccd1 _9302_/X sky130_fd_sc_hd__mux2_1
X_9233_ _9232_/X _7786_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9233_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7494_ _7494_/A _7494_/B vssd1 vssd1 vccd1 vccd1 _7494_/X sky130_fd_sc_hd__or2_1
XFILLER_173_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6445_ _6339_/Y _6443_/Y _6376_/B vssd1 vssd1 vccd1 vccd1 _6447_/A sky130_fd_sc_hd__o21ai_1
X_9164_ _6273_/X input33/X _9170_/S vssd1 vssd1 vccd1 vccd1 _9164_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6376_ _9758_/Q _6376_/B vssd1 vssd1 vccd1 vccd1 _6377_/B sky130_fd_sc_hd__or2_2
X_8115_ _9541_/Q _8069_/B _8070_/B vssd1 vssd1 vccd1 vccd1 _8115_/X sky130_fd_sc_hd__a21bo_1
X_9095_ _6564_/X _6566_/Y _9683_/Q vssd1 vssd1 vccd1 vccd1 _9095_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5327_ _5327_/A _5388_/A vssd1 vssd1 vccd1 vccd1 _5384_/A sky130_fd_sc_hd__or2_1
X_8046_ _8046_/A _8046_/B vssd1 vssd1 vccd1 vccd1 _8046_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5258_ _5258_/A _5258_/B vssd1 vssd1 vccd1 vccd1 _9746_/D sky130_fd_sc_hd__nor2_1
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5189_ _9763_/Q _5203_/A input22/X _5205_/A _5187_/X vssd1 vssd1 vccd1 vccd1 _9763_/D
+ sky130_fd_sc_hd__o221a_1
X_8948_ _8941_/X _8947_/X _8941_/X _8947_/X vssd1 vssd1 vccd1 vccd1 _8948_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8879_ _8874_/X _8878_/X _8874_/X _8878_/X vssd1 vssd1 vccd1 vccd1 _8881_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6230_ _9581_/Q vssd1 vssd1 vccd1 vccd1 _8017_/A sky130_fd_sc_hd__inv_2
X_6161_ _6152_/X _6155_/X _6160_/X vssd1 vssd1 vccd1 vccd1 _6161_/Y sky130_fd_sc_hd__o21ai_2
X_5112_ _9797_/Q vssd1 vssd1 vccd1 vccd1 _5112_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6092_ _7999_/A _9648_/Q vssd1 vssd1 vccd1 vccd1 _6095_/A sky130_fd_sc_hd__nor2_1
X_9920_ _9923_/CLK _9920_/D vssd1 vssd1 vccd1 vccd1 _9920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5043_ _5214_/A vssd1 vssd1 vccd1 vccd1 _5070_/A sky130_fd_sc_hd__buf_6
XFILLER_38_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9851_ _9858_/CLK _9851_/D vssd1 vssd1 vccd1 vccd1 _9851_/Q sky130_fd_sc_hd__dfxtp_2
X_8802_ _8800_/A _8725_/B _5843_/X _8610_/B vssd1 vssd1 vccd1 vccd1 _8803_/A sky130_fd_sc_hd__o211a_1
XFILLER_80_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9782_ _9819_/CLK _9782_/D vssd1 vssd1 vccd1 vccd1 _9782_/Q sky130_fd_sc_hd__dfxtp_1
X_6994_ _6969_/A _6971_/B _7006_/A _7005_/B vssd1 vssd1 vccd1 vccd1 _6995_/B sky130_fd_sc_hd__o22a_1
XFILLER_92_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8733_ _8821_/A _8875_/D vssd1 vssd1 vccd1 vccd1 _8823_/C sky130_fd_sc_hd__or2_2
XFILLER_80_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5945_ _5959_/A vssd1 vssd1 vccd1 vccd1 _5945_/X sky130_fd_sc_hd__clkbuf_2
X_8664_ _8662_/Y _8663_/Y _8662_/Y _8663_/Y vssd1 vssd1 vccd1 vccd1 _8709_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_178_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5876_ _9621_/Q _5865_/A _4860_/A _5866_/A _5875_/X vssd1 vssd1 vccd1 vccd1 _9621_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_40_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4827_ _9262_/X _4822_/X _9906_/Q _4824_/X _4817_/X vssd1 vssd1 vccd1 vccd1 _9906_/D
+ sky130_fd_sc_hd__o221a_1
X_7615_ _7600_/A _7600_/B _7601_/B vssd1 vssd1 vccd1 vccd1 _7615_/X sky130_fd_sc_hd__a21bo_1
X_8595_ _8542_/X _8550_/Y _8551_/X _8552_/X vssd1 vssd1 vccd1 vccd1 _8596_/B sky130_fd_sc_hd__o22a_4
XFILLER_178_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4758_ _5891_/A vssd1 vssd1 vccd1 vccd1 _5916_/A sky130_fd_sc_hd__buf_4
XFILLER_119_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7546_ _7543_/X _7545_/X _7543_/X _7545_/X vssd1 vssd1 vccd1 vccd1 _7546_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_181_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7477_ _7477_/A _7477_/B vssd1 vssd1 vccd1 vccd1 _7537_/B sky130_fd_sc_hd__or2_1
XFILLER_161_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9216_ _9821_/Q _7647_/Y _9528_/Q vssd1 vssd1 vccd1 vccd1 _9216_/X sky130_fd_sc_hd__mux2_1
X_6428_ _6428_/A vssd1 vssd1 vccd1 vccd1 _6535_/B sky130_fd_sc_hd__inv_2
XFILLER_134_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9147_ _6180_/Y input46/X _9148_/S vssd1 vssd1 vccd1 vccd1 _9147_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6359_ _8051_/A _9752_/Q vssd1 vssd1 vccd1 vccd1 _6359_/Y sky130_fd_sc_hd__nor2_1
X_9078_ _9077_/X _7833_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9078_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8029_ _8029_/A _8033_/B vssd1 vssd1 vccd1 vccd1 _8029_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5730_ _9676_/Q _9659_/Q _6582_/A _5729_/Y vssd1 vssd1 vccd1 vccd1 _5730_/X sky130_fd_sc_hd__a22o_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5661_ _9689_/Q _5658_/X _6556_/A _5650_/X _5660_/X vssd1 vssd1 vccd1 vccd1 _9689_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7400_ _7400_/A _7400_/B _7400_/C vssd1 vssd1 vccd1 vccd1 _7400_/X sky130_fd_sc_hd__or3_1
XFILLER_175_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5592_ _5494_/X _5532_/X _5494_/X _5532_/X vssd1 vssd1 vccd1 vccd1 _5592_/Y sky130_fd_sc_hd__a2bb2oi_2
X_8380_ _9697_/Q vssd1 vssd1 vccd1 vccd1 _8381_/A sky130_fd_sc_hd__inv_2
XFILLER_190_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7331_ _7331_/A _7400_/B _7331_/C vssd1 vssd1 vccd1 vccd1 _7331_/X sky130_fd_sc_hd__or3_1
XFILLER_209_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7262_ _7256_/A _7428_/A _7255_/Y _7253_/A _7261_/Y vssd1 vssd1 vccd1 vccd1 _7262_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_143_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9001_ _5112_/Y _7723_/X _9480_/S vssd1 vssd1 vccd1 vccd1 _9001_/X sky130_fd_sc_hd__mux2_1
X_6213_ _6221_/A _6221_/B _6204_/Y _6212_/X vssd1 vssd1 vccd1 vccd1 _6213_/X sky130_fd_sc_hd__o31a_1
X_7193_ _7187_/A _7503_/A _7186_/Y _7184_/A _7192_/Y vssd1 vssd1 vccd1 vccd1 _7193_/X
+ sky130_fd_sc_hd__o32a_1
X_6144_ _6125_/Y _6143_/X _6150_/A vssd1 vssd1 vccd1 vccd1 _6144_/Y sky130_fd_sc_hd__o21ai_1
XINSDIODE2_16 input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6075_ _9859_/Q _6074_/B _6074_/Y vssd1 vssd1 vccd1 vccd1 _6076_/A sky130_fd_sc_hd__a21oi_4
X_9903_ _9903_/CLK _9903_/D vssd1 vssd1 vccd1 vccd1 _9903_/Q sky130_fd_sc_hd__dfxtp_1
X_5026_ _5026_/A vssd1 vssd1 vccd1 vccd1 _5026_/X sky130_fd_sc_hd__buf_4
X_9834_ _9923_/CLK _9834_/D vssd1 vssd1 vccd1 vccd1 _9834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6977_ _6973_/X _6976_/Y _6973_/X _6976_/Y vssd1 vssd1 vccd1 vccd1 _6977_/X sky130_fd_sc_hd__a2bb2o_1
X_9765_ _9916_/CLK _9765_/D vssd1 vssd1 vccd1 vccd1 _9765_/Q sky130_fd_sc_hd__dfxtp_2
X_5928_ _9167_/X _5921_/X _9591_/Q _5924_/X vssd1 vssd1 vccd1 vccd1 _9591_/D sky130_fd_sc_hd__a22o_1
XFILLER_179_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8716_ _8633_/A _8714_/Y _8677_/Y _8674_/Y _8715_/X vssd1 vssd1 vccd1 vccd1 _8717_/A
+ sky130_fd_sc_hd__a32o_1
X_9696_ _9699_/CLK _9696_/D vssd1 vssd1 vccd1 vccd1 _9696_/Q sky130_fd_sc_hd__dfxtp_1
X_5859_ _5858_/X _5847_/A _5039_/X _5848_/A _5853_/X vssd1 vssd1 vccd1 vccd1 _9628_/D
+ sky130_fd_sc_hd__o221a_1
X_8647_ _9693_/Q _8386_/B _8386_/Y vssd1 vssd1 vccd1 vccd1 _8647_/X sky130_fd_sc_hd__a21o_1
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8578_ _8574_/X _8577_/X _8574_/X _8577_/X vssd1 vssd1 vccd1 vccd1 _8578_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7529_ _7527_/X _7528_/X _7527_/X _7528_/X vssd1 vssd1 vccd1 vccd1 _7529_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_181_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7880_ _4786_/X _7679_/B _7879_/Y vssd1 vssd1 vccd1 vccd1 _7880_/X sky130_fd_sc_hd__a21o_1
X_6900_ _6888_/A _6888_/B _6925_/A vssd1 vssd1 vccd1 vccd1 _6903_/A sky130_fd_sc_hd__a21o_1
X_6831_ _6819_/A _6819_/B _6846_/A vssd1 vssd1 vccd1 vccd1 _6834_/A sky130_fd_sc_hd__a21o_1
X_9550_ _9923_/CLK _9550_/D vssd1 vssd1 vccd1 vccd1 _9550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8501_ _8576_/C vssd1 vssd1 vccd1 vccd1 _8529_/C sky130_fd_sc_hd__inv_2
X_6762_ _6749_/X _6750_/X _6749_/X _6750_/X vssd1 vssd1 vccd1 vccd1 _6762_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9481_ _9480_/X _6348_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _9481_/X sky130_fd_sc_hd__mux2_1
X_5713_ _9665_/Q vssd1 vssd1 vccd1 vccd1 _5713_/Y sky130_fd_sc_hd__inv_2
X_6693_ _6760_/B vssd1 vssd1 vccd1 vccd1 _6766_/B sky130_fd_sc_hd__clkbuf_2
X_8432_ _8432_/A _8432_/B vssd1 vssd1 vccd1 vccd1 _8446_/A sky130_fd_sc_hd__or2_1
X_5644_ _5644_/A vssd1 vssd1 vccd1 vccd1 _5689_/A sky130_fd_sc_hd__clkbuf_2
X_8363_ _8363_/A _8363_/B _8361_/X _8362_/X vssd1 vssd1 vccd1 vccd1 _8375_/C sky130_fd_sc_hd__or4bb_4
XFILLER_163_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5575_ _9710_/Q vssd1 vssd1 vccd1 vccd1 _7648_/A sky130_fd_sc_hd__inv_2
X_7314_ _7314_/A _9473_/X vssd1 vssd1 vccd1 vccd1 _7314_/X sky130_fd_sc_hd__or2_1
XFILLER_191_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8294_ _7885_/X _8207_/X _7892_/A _8206_/X _8293_/X vssd1 vssd1 vccd1 vccd1 _8294_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_131_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7245_ _7245_/A _7245_/B vssd1 vssd1 vccd1 vccd1 _7256_/A sky130_fd_sc_hd__or2_1
X_7176_ _7176_/A _7176_/B vssd1 vssd1 vccd1 vccd1 _7187_/A sky130_fd_sc_hd__or2_2
XFILLER_98_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6127_ _6146_/A vssd1 vssd1 vccd1 vccd1 _6148_/A sky130_fd_sc_hd__inv_2
XFILLER_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6058_ _9856_/Q _6041_/Y _6049_/A vssd1 vssd1 vccd1 vccd1 _6059_/A sky130_fd_sc_hd__o21ai_2
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5009_ _9830_/Q _5003_/X input25/X _5004_/X _5008_/X vssd1 vssd1 vccd1 vccd1 _9830_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_199_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9817_ _9819_/CLK _9817_/D vssd1 vssd1 vccd1 vccd1 _9817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9748_ _9750_/CLK _9748_/D vssd1 vssd1 vccd1 vccd1 _9748_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_121_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9679_ _9699_/CLK _9679_/D vssd1 vssd1 vccd1 vccd1 _9679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_31_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _9861_/CLK sky130_fd_sc_hd__clkbuf_16
X_5360_ _5360_/A vssd1 vssd1 vccd1 vccd1 _9727_/D sky130_fd_sc_hd__inv_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5291_ _9738_/Q _5291_/B vssd1 vssd1 vccd1 vccd1 _5291_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7030_ _7030_/A _7030_/B vssd1 vssd1 vccd1 vccd1 _7030_/X sky130_fd_sc_hd__or2_1
XFILLER_141_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8981_ _7981_/X _6055_/B _9504_/S vssd1 vssd1 vccd1 vccd1 _8981_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7932_ _8471_/A vssd1 vssd1 vccd1 vccd1 _8534_/A sky130_fd_sc_hd__buf_1
XFILLER_95_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7863_ _7863_/A vssd1 vssd1 vccd1 vccd1 _7863_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7794_ _8324_/A _7789_/Y _7797_/B _7785_/X vssd1 vssd1 vccd1 vccd1 _7794_/X sky130_fd_sc_hd__o211a_1
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9602_ _9895_/CLK _9602_/D vssd1 vssd1 vccd1 vccd1 _9602_/Q sky130_fd_sc_hd__dfxtp_1
X_6814_ _6814_/A _6883_/B _6814_/C vssd1 vssd1 vccd1 vccd1 _6814_/X sky130_fd_sc_hd__or3_1
XFILLER_211_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9533_ _9796_/CLK _9533_/D vssd1 vssd1 vccd1 vccd1 _9533_/Q sky130_fd_sc_hd__dfxtp_1
X_6745_ _6739_/A _6911_/A _6738_/Y _6736_/A _6744_/Y vssd1 vssd1 vccd1 vccd1 _6745_/X
+ sky130_fd_sc_hd__o32a_1
XPHY_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9464_ _6582_/X _6584_/Y _9683_/Q vssd1 vssd1 vccd1 vccd1 _9464_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6676_ _6654_/X _6675_/X _6654_/X _6675_/X vssd1 vssd1 vccd1 vccd1 _6676_/X sky130_fd_sc_hd__a2bb2o_1
X_8415_ _5515_/X _6573_/X _8396_/X _8397_/Y vssd1 vssd1 vccd1 vccd1 _8415_/X sky130_fd_sc_hd__a31o_1
XFILLER_109_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5627_ _5627_/A _8436_/C vssd1 vssd1 vccd1 vccd1 _5627_/X sky130_fd_sc_hd__and2_1
X_9395_ _8700_/X _8698_/A _9477_/S vssd1 vssd1 vccd1 vccd1 _9395_/X sky130_fd_sc_hd__mux2_1
X_8346_ _8346_/A _8346_/B _8344_/X _8345_/X vssd1 vssd1 vccd1 vccd1 _8375_/D sky130_fd_sc_hd__or4bb_4
XFILLER_117_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5558_ _5553_/X _5554_/Y _5555_/Y _7652_/A _5557_/X vssd1 vssd1 vccd1 vccd1 _5559_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_144_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8277_ _7835_/A _8230_/X _8276_/Y vssd1 vssd1 vccd1 vccd1 _8277_/X sky130_fd_sc_hd__a21o_1
XFILLER_116_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7228_ _7273_/B vssd1 vssd1 vccd1 vccd1 _7291_/B sky130_fd_sc_hd__clkbuf_2
X_5489_ _5420_/X _5457_/X _5420_/X _5457_/X vssd1 vssd1 vccd1 vccd1 _5489_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7159_ _9430_/X vssd1 vssd1 vccd1 vccd1 _7210_/B sky130_fd_sc_hd__inv_2
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4860_ _4860_/A vssd1 vssd1 vccd1 vccd1 _4860_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_177_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4791_ _4830_/A vssd1 vssd1 vccd1 vccd1 _4791_/X sky130_fd_sc_hd__clkbuf_2
X_6530_ _6550_/A vssd1 vssd1 vccd1 vccd1 _6535_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6461_ _9789_/Q _6525_/B _9788_/Q _6522_/B _6446_/X vssd1 vssd1 vccd1 vccd1 _6462_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_9_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6392_ _9774_/Q _6407_/A vssd1 vssd1 vccd1 vccd1 _6393_/B sky130_fd_sc_hd__or2_2
X_8200_ _8200_/A _8200_/B vssd1 vssd1 vccd1 vccd1 _8200_/Y sky130_fd_sc_hd__nor2_1
X_9180_ _6519_/Y _9785_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9534_/D sky130_fd_sc_hd__mux2_1
X_5412_ _5412_/A _5412_/B vssd1 vssd1 vccd1 vccd1 _5412_/Y sky130_fd_sc_hd__nor2_1
X_8131_ _8134_/B vssd1 vssd1 vccd1 vccd1 _8131_/Y sky130_fd_sc_hd__inv_2
X_5343_ _5343_/A vssd1 vssd1 vccd1 vccd1 _9731_/D sky130_fd_sc_hd__inv_2
X_8062_ _9534_/Q _8062_/B vssd1 vssd1 vccd1 vccd1 _8063_/B sky130_fd_sc_hd__or2_1
XFILLER_102_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5274_ _9896_/Q vssd1 vssd1 vccd1 vccd1 _5275_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7013_ _6964_/A _6964_/B _6964_/X vssd1 vssd1 vccd1 vccd1 _7013_/X sky130_fd_sc_hd__a21bo_1
XFILLER_83_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8964_ _8950_/Y _8963_/Y _8950_/Y _8963_/Y vssd1 vssd1 vccd1 vccd1 _8964_/X sky130_fd_sc_hd__a2bb2o_2
X_8895_ _8895_/A _8895_/B vssd1 vssd1 vccd1 vccd1 _8895_/X sky130_fd_sc_hd__or2_1
XFILLER_102_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7915_ input3/X input6/X _5881_/A _8008_/B _5709_/B vssd1 vssd1 vccd1 vccd1 _7991_/A
+ sky130_fd_sc_hd__o311a_2
X_7846_ _7846_/A vssd1 vssd1 vccd1 vccd1 _7846_/Y sky130_fd_sc_hd__inv_2
XPHY_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4989_ _9842_/Q _4985_/X input39/X _4987_/X _4974_/X vssd1 vssd1 vccd1 vccd1 _9842_/D
+ sky130_fd_sc_hd__o221a_1
X_7777_ _7777_/A vssd1 vssd1 vccd1 vccd1 _7779_/A sky130_fd_sc_hd__inv_2
XPHY_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9516_ _9634_/CLK input1/X vssd1 vssd1 vccd1 vccd1 _9517_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_184_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6728_ _6728_/A _6728_/B vssd1 vssd1 vccd1 vccd1 _6739_/A sky130_fd_sc_hd__or2_1
XPHY_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9447_ _9811_/Q _9928_/Q _9480_/S vssd1 vssd1 vccd1 vccd1 _9447_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6659_ _6646_/X _6647_/X _6646_/X _6647_/X vssd1 vssd1 vccd1 vccd1 _6659_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9378_ _8447_/Y _8444_/X _9477_/S vssd1 vssd1 vccd1 vccd1 _9378_/X sky130_fd_sc_hd__mux2_4
XFILLER_137_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8329_ _7769_/Y _9537_/Q _7715_/X _9544_/Q vssd1 vssd1 vccd1 vccd1 _8331_/B sky130_fd_sc_hd__a22o_1
XFILLER_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput37 io_wb_dat_i[29] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__buf_4
XFILLER_167_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput26 io_wb_dat_i[19] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_4
XPHY_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput15 io_wb_cs_i vssd1 vssd1 vccd1 vccd1 _4855_/B sky130_fd_sc_hd__buf_2
XFILLER_128_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput48 io_wb_we_i vssd1 vssd1 vccd1 vccd1 _4744_/A sky130_fd_sc_hd__buf_2
XFILLER_143_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5961_ _9145_/X _5958_/X _9568_/Q _5959_/X vssd1 vssd1 vccd1 vccd1 _9568_/D sky130_fd_sc_hd__a22o_1
XFILLER_206_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8680_ _8655_/X _8679_/X _8655_/X _8679_/X vssd1 vssd1 vccd1 vccd1 _8680_/X sky130_fd_sc_hd__a2bb2o_1
X_7700_ _7891_/A _5162_/X _4816_/X _6333_/Y vssd1 vssd1 vccd1 vccd1 _7700_/X sky130_fd_sc_hd__o22a_1
XFILLER_80_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4912_ _5662_/A vssd1 vssd1 vccd1 vccd1 _4912_/X sky130_fd_sc_hd__clkbuf_2
X_5892_ _5890_/X _5884_/X _4978_/A _5885_/X _5891_/X vssd1 vssd1 vccd1 vccd1 _9615_/D
+ sky130_fd_sc_hd__o221a_1
X_7631_ _7592_/A _7592_/B _7593_/B vssd1 vssd1 vccd1 vccd1 _7631_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_178_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4843_ _7657_/A vssd1 vssd1 vccd1 vccd1 _4843_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4774_ _9925_/Q vssd1 vssd1 vccd1 vccd1 _7682_/A sky130_fd_sc_hd__buf_2
XFILLER_166_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7562_ _7553_/A _7553_/B _7553_/Y vssd1 vssd1 vccd1 vccd1 _7562_/Y sky130_fd_sc_hd__o21ai_1
X_6513_ _9807_/Q _6546_/B _9806_/Q _6545_/B _6512_/Y vssd1 vssd1 vccd1 vccd1 _6513_/X
+ sky130_fd_sc_hd__o221a_1
X_9301_ _9300_/X _7870_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9301_/X sky130_fd_sc_hd__mux2_1
X_7493_ _7491_/X _7492_/X _7491_/X _7492_/X vssd1 vssd1 vccd1 vccd1 _7493_/Y sky130_fd_sc_hd__a2bb2oi_1
X_9232_ _9750_/Q _9231_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9232_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6444_ _6341_/A _6374_/B _6443_/Y vssd1 vssd1 vccd1 vccd1 _6522_/B sky130_fd_sc_hd__a21oi_2
XFILLER_9_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9163_ _6269_/Y input32/X _9170_/S vssd1 vssd1 vccd1 vccd1 _9163_/X sky130_fd_sc_hd__mux2_1
X_6375_ _9757_/Q _6443_/A vssd1 vssd1 vccd1 vccd1 _6376_/B sky130_fd_sc_hd__or2_1
XFILLER_161_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8114_ _9542_/Q _8070_/B _8112_/Y vssd1 vssd1 vccd1 vccd1 _8114_/X sky130_fd_sc_hd__a21o_1
X_9094_ _8391_/B _6563_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9094_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5326_ _9719_/Q _5392_/B vssd1 vssd1 vccd1 vccd1 _5388_/A sky130_fd_sc_hd__nand2_1
X_8045_ _9479_/X _8045_/B vssd1 vssd1 vccd1 vccd1 _8045_/Y sky130_fd_sc_hd__nor2_1
X_5257_ _5251_/B _5253_/Y _9746_/Q vssd1 vssd1 vccd1 vccd1 _5258_/B sky130_fd_sc_hd__a21oi_1
XFILLER_102_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5188_ _6353_/A _5178_/X input23/X _5179_/X _5187_/X vssd1 vssd1 vccd1 vccd1 _9764_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_87_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8947_ _8942_/Y _8946_/X _8942_/Y _8946_/X vssd1 vssd1 vccd1 vccd1 _8947_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8878_ _8878_/A _8878_/B vssd1 vssd1 vccd1 vccd1 _8878_/X sky130_fd_sc_hd__or2_1
XPHY_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7829_ _7829_/A vssd1 vssd1 vccd1 vccd1 _7829_/Y sky130_fd_sc_hd__inv_2
XPHY_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6160_ _7949_/A _6135_/A _7957_/A _6135_/A vssd1 vssd1 vccd1 vccd1 _6160_/X sky130_fd_sc_hd__o22a_1
X_5111_ _5115_/A _5111_/B vssd1 vssd1 vccd1 vccd1 _9798_/D sky130_fd_sc_hd__nor2_1
X_6091_ _9861_/Q vssd1 vssd1 vccd1 vccd1 _7999_/A sky130_fd_sc_hd__inv_2
X_5042_ _9812_/Q _5003_/A _5041_/X _5004_/A _5036_/X vssd1 vssd1 vccd1 vccd1 _9812_/D
+ sky130_fd_sc_hd__o221a_1
X_9850_ _9858_/CLK _9850_/D vssd1 vssd1 vccd1 vccd1 _9850_/Q sky130_fd_sc_hd__dfxtp_2
X_8801_ _8801_/A vssd1 vssd1 vccd1 vccd1 _8893_/C sky130_fd_sc_hd__inv_2
XFILLER_198_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9781_ _9819_/CLK _9781_/D vssd1 vssd1 vccd1 vccd1 _9781_/Q sky130_fd_sc_hd__dfxtp_1
X_6993_ _6990_/X _6992_/X _6990_/X _6992_/X vssd1 vssd1 vccd1 vccd1 _6993_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8732_ _8730_/X _8731_/X _8730_/X _8731_/X vssd1 vssd1 vccd1 vccd1 _8732_/X sky130_fd_sc_hd__a2bb2o_1
X_5944_ _5958_/A vssd1 vssd1 vccd1 vccd1 _5944_/X sky130_fd_sc_hd__clkbuf_2
X_8663_ _8609_/A _8611_/Y _8612_/X _8617_/X vssd1 vssd1 vccd1 vccd1 _8663_/Y sky130_fd_sc_hd__o22ai_2
X_5875_ _5891_/A vssd1 vssd1 vccd1 vccd1 _5875_/X sky130_fd_sc_hd__clkbuf_2
X_8594_ _8593_/A _8593_/B _8593_/Y vssd1 vssd1 vccd1 vccd1 _8596_/A sky130_fd_sc_hd__a21o_2
XFILLER_166_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4826_ _9266_/X _4822_/X _9907_/Q _4824_/X _4817_/X vssd1 vssd1 vccd1 vccd1 _9907_/D
+ sky130_fd_sc_hd__o221a_1
X_7614_ _7077_/A _7077_/B _7078_/B vssd1 vssd1 vccd1 vccd1 _7614_/X sky130_fd_sc_hd__a21bo_1
XFILLER_61_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7545_ _7492_/C _7210_/B _7273_/A _7135_/Y _7544_/X vssd1 vssd1 vccd1 vccd1 _7545_/X
+ sky130_fd_sc_hd__a41o_1
X_4757_ _5790_/A vssd1 vssd1 vccd1 vccd1 _5891_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7476_ _7438_/X _7448_/X _7474_/X _7475_/X vssd1 vssd1 vccd1 vccd1 _7476_/X sky130_fd_sc_hd__o22a_1
X_9215_ _9820_/Q _7646_/Y _9528_/Q vssd1 vssd1 vccd1 vccd1 _9215_/X sky130_fd_sc_hd__mux2_1
X_6427_ _6427_/A vssd1 vssd1 vccd1 vccd1 _6534_/B sky130_fd_sc_hd__inv_2
X_6358_ _8183_/A vssd1 vssd1 vccd1 vccd1 _8051_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_122_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9146_ _6173_/X _5026_/A _9155_/S vssd1 vssd1 vccd1 vccd1 _9146_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5309_ _5305_/Y _5224_/A _5308_/Y _5275_/A _5238_/A vssd1 vssd1 vccd1 vccd1 _5310_/A
+ sky130_fd_sc_hd__o32a_1
X_6289_ _6288_/A _6288_/B _6296_/A vssd1 vssd1 vccd1 vccd1 _6289_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_102_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9077_ _9761_/Q _9076_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9077_/X sky130_fd_sc_hd__mux2_1
X_8028_ _9481_/X _8037_/B vssd1 vssd1 vccd1 vccd1 _8028_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5660_ _5660_/A vssd1 vssd1 vccd1 vccd1 _5660_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5591_ _5609_/A _5591_/B vssd1 vssd1 vccd1 vccd1 _9708_/D sky130_fd_sc_hd__nor2_1
XFILLER_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7330_ _7330_/A vssd1 vssd1 vccd1 vccd1 _7331_/C sky130_fd_sc_hd__inv_2
XFILLER_116_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7261_ _7261_/A _7427_/B vssd1 vssd1 vccd1 vccd1 _7261_/Y sky130_fd_sc_hd__nor2_1
XFILLER_209_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9000_ _8999_/X _9523_/Q _9155_/S vssd1 vssd1 vccd1 vccd1 _9000_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6212_ _7997_/A _6201_/X _8001_/A _6201_/X vssd1 vssd1 vccd1 vccd1 _6212_/X sky130_fd_sc_hd__o22a_1
XFILLER_131_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7192_ _7192_/A _7502_/B vssd1 vssd1 vccd1 vccd1 _7192_/Y sky130_fd_sc_hd__nor2_1
X_6143_ _6193_/A vssd1 vssd1 vccd1 vccd1 _6143_/X sky130_fd_sc_hd__buf_6
XFILLER_124_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6074_ _9859_/Q _6074_/B vssd1 vssd1 vccd1 vccd1 _6074_/Y sky130_fd_sc_hd__nor2_2
XINSDIODE2_17 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9902_ _9903_/CLK _9902_/D vssd1 vssd1 vccd1 vccd1 _9902_/Q sky130_fd_sc_hd__dfxtp_2
X_5025_ _9820_/Q _5019_/X input46/X _5020_/X _5024_/X vssd1 vssd1 vccd1 vccd1 _9820_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9833_ _9833_/CLK _9833_/D vssd1 vssd1 vccd1 vccd1 _9833_/Q sky130_fd_sc_hd__dfxtp_1
X_6976_ _6974_/Y _6975_/X _6974_/Y _6975_/X vssd1 vssd1 vccd1 vccd1 _6976_/Y sky130_fd_sc_hd__o2bb2ai_1
X_9764_ _9916_/CLK _9764_/D vssd1 vssd1 vccd1 vccd1 _9764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5927_ _9168_/X _5921_/X _9592_/Q _5924_/X vssd1 vssd1 vccd1 vccd1 _9592_/D sky130_fd_sc_hd__a22o_1
X_8715_ _8715_/A _8715_/B vssd1 vssd1 vccd1 vccd1 _8715_/X sky130_fd_sc_hd__or2_1
X_9695_ _9699_/CLK _9695_/D vssd1 vssd1 vccd1 vccd1 _9695_/Q sky130_fd_sc_hd__dfxtp_1
X_5858_ _9628_/Q vssd1 vssd1 vccd1 vccd1 _5858_/X sky130_fd_sc_hd__buf_2
XFILLER_166_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8646_ _8645_/A _8645_/B _8695_/A vssd1 vssd1 vccd1 vccd1 _8646_/X sky130_fd_sc_hd__a21bo_1
XFILLER_70_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8577_ _8528_/X _8529_/X _8530_/X _8532_/X _8576_/X vssd1 vssd1 vccd1 vccd1 _8577_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_186_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5789_ _5749_/X _5788_/X _5749_/X _5788_/X vssd1 vssd1 vccd1 vccd1 _7089_/A sky130_fd_sc_hd__o2bb2a_2
X_4809_ _4834_/A vssd1 vssd1 vccd1 vccd1 _4809_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7528_ _7509_/X _7514_/X _7509_/X _7514_/X vssd1 vssd1 vccd1 vccd1 _7528_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7459_ _7419_/A _7419_/B _7420_/B vssd1 vssd1 vccd1 vccd1 _7459_/X sky130_fd_sc_hd__a21bo_1
XFILLER_162_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9129_ _9866_/Q _9882_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9129_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6830_ _6830_/A vssd1 vssd1 vccd1 vccd1 _6846_/A sky130_fd_sc_hd__inv_2
XFILLER_211_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6761_ _6751_/X _6752_/X _6759_/X _6760_/X vssd1 vssd1 vccd1 vccd1 _6761_/X sky130_fd_sc_hd__o22a_1
XFILLER_35_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8500_ _9378_/X vssd1 vssd1 vccd1 vccd1 _8500_/Y sky130_fd_sc_hd__inv_2
X_5712_ _9682_/Q vssd1 vssd1 vccd1 vccd1 _6598_/A sky130_fd_sc_hd__inv_2
XFILLER_203_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9480_ _6318_/B _7869_/A _9480_/S vssd1 vssd1 vccd1 vccd1 _9480_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6692_ _9092_/X vssd1 vssd1 vccd1 vccd1 _6760_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_8431_ _8432_/B vssd1 vssd1 vccd1 vccd1 _8431_/Y sky130_fd_sc_hd__inv_2
X_5643_ _9695_/Q _5631_/X _6578_/A _5635_/X _5632_/X vssd1 vssd1 vccd1 vccd1 _9695_/D
+ sky130_fd_sc_hd__o221a_1
X_8362_ _9926_/Q _8092_/Y _7684_/A _8048_/Y vssd1 vssd1 vccd1 vccd1 _8362_/X sky130_fd_sc_hd__o22a_1
XFILLER_148_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5574_ _5574_/A _5574_/B vssd1 vssd1 vccd1 vccd1 _5574_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7313_ _7334_/A _9475_/X _7313_/C _7334_/B vssd1 vssd1 vccd1 vccd1 _7313_/X sky130_fd_sc_hd__or4_4
X_8293_ _7887_/A _8207_/X _7881_/X _8208_/Y _8292_/X vssd1 vssd1 vccd1 vccd1 _8293_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7244_ _7233_/A _7233_/B _7233_/X vssd1 vssd1 vccd1 vccd1 _7245_/B sky130_fd_sc_hd__a21bo_1
XFILLER_104_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7175_ _7164_/A _7164_/B _7164_/X vssd1 vssd1 vccd1 vccd1 _7176_/B sky130_fd_sc_hd__a21bo_1
XFILLER_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6126_ _6126_/A vssd1 vssd1 vccd1 vccd1 _6146_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6057_ _6057_/A vssd1 vssd1 vccd1 vccd1 _6057_/Y sky130_fd_sc_hd__inv_2
X_5008_ _5036_/A vssd1 vssd1 vccd1 vccd1 _5008_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9816_ _9819_/CLK _9816_/D vssd1 vssd1 vccd1 vccd1 _9816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9747_ _9887_/CLK _9747_/D vssd1 vssd1 vccd1 vccd1 _9747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6959_ _6921_/X _6931_/X _6932_/X _6958_/X vssd1 vssd1 vccd1 vccd1 _6959_/X sky130_fd_sc_hd__o22a_1
XFILLER_53_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9678_ _9699_/CLK _9678_/D vssd1 vssd1 vccd1 vccd1 _9678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8629_ _8629_/A vssd1 vssd1 vccd1 vccd1 _8629_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5290_ _5290_/A vssd1 vssd1 vccd1 vccd1 _5291_/B sky130_fd_sc_hd__inv_2
XFILLER_99_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8980_ _8979_/X _6341_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _8980_/X sky130_fd_sc_hd__mux2_2
XFILLER_121_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7931_ _9629_/Q vssd1 vssd1 vccd1 vccd1 _8471_/A sky130_fd_sc_hd__inv_2
XFILLER_82_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7862_ _4802_/X _7857_/Y _7860_/X _7865_/B vssd1 vssd1 vccd1 vccd1 _7862_/X sky130_fd_sc_hd__o211a_1
X_9601_ _9895_/CLK _9601_/D vssd1 vssd1 vccd1 vccd1 _9601_/Q sky130_fd_sc_hd__dfxtp_1
X_7793_ _7793_/A _7793_/B vssd1 vssd1 vccd1 vccd1 _7797_/B sky130_fd_sc_hd__or2_2
X_6813_ _6813_/A vssd1 vssd1 vccd1 vccd1 _6814_/C sky130_fd_sc_hd__inv_2
XFILLER_211_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9532_ _9796_/CLK _9532_/D vssd1 vssd1 vccd1 vccd1 _9532_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6744_ _6744_/A _6910_/B vssd1 vssd1 vccd1 vccd1 _6744_/Y sky130_fd_sc_hd__nor2_1
XFILLER_195_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6675_ _6669_/A _6992_/A _6668_/Y _6666_/A _6674_/Y vssd1 vssd1 vccd1 vccd1 _6675_/X
+ sky130_fd_sc_hd__o32a_1
X_9463_ _8386_/B _6583_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9463_/X sky130_fd_sc_hd__mux2_2
XFILLER_50_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5626_ _5626_/A vssd1 vssd1 vccd1 vccd1 _5626_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8414_ _8411_/X _8413_/X _8411_/X _8413_/X vssd1 vssd1 vccd1 vccd1 _9490_/S sky130_fd_sc_hd__o2bb2ai_4
XFILLER_136_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9394_ _8794_/X _8792_/A _9490_/S vssd1 vssd1 vccd1 vccd1 _9394_/X sky130_fd_sc_hd__mux2_1
X_8345_ _4798_/X _8102_/Y _4794_/X _8334_/Y vssd1 vssd1 vccd1 vccd1 _8345_/X sky130_fd_sc_hd__o22a_1
XFILLER_117_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5557_ _5644_/A vssd1 vssd1 vccd1 vccd1 _5557_/X sky130_fd_sc_hd__buf_2
XFILLER_132_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5488_ _9385_/X _5487_/X _9385_/X _5487_/X vssd1 vssd1 vccd1 vccd1 _5582_/A sky130_fd_sc_hd__a2bb2oi_1
XFILLER_104_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8276_ _9910_/Q _8233_/Y _8275_/X vssd1 vssd1 vccd1 vccd1 _8276_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7227_ _9471_/X vssd1 vssd1 vccd1 vccd1 _7273_/B sky130_fd_sc_hd__inv_2
XFILLER_116_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7158_ _7195_/A _9424_/X vssd1 vssd1 vccd1 vccd1 _7165_/C sky130_fd_sc_hd__nor2_1
XFILLER_86_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6109_ _9863_/Q vssd1 vssd1 vccd1 vccd1 _8008_/A sky130_fd_sc_hd__inv_2
X_7089_ _7089_/A _7089_/B vssd1 vssd1 vccd1 vccd1 _7107_/B sky130_fd_sc_hd__or2_2
XFILLER_132_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4790_ _9920_/Q vssd1 vssd1 vccd1 vccd1 _4790_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6460_ _6465_/C _6465_/B _6458_/Y _6463_/C vssd1 vssd1 vccd1 vccd1 _6460_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6391_ _9773_/Q _8203_/A vssd1 vssd1 vccd1 vccd1 _6407_/A sky130_fd_sc_hd__or2_1
X_5411_ _9346_/X vssd1 vssd1 vccd1 vccd1 _5412_/B sky130_fd_sc_hd__inv_2
X_8130_ _8058_/Y _8129_/X _8058_/Y _8129_/X vssd1 vssd1 vccd1 vccd1 _8134_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_126_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5342_ _9731_/Q _5313_/X _5340_/C _5338_/Y _5341_/Y vssd1 vssd1 vccd1 vccd1 _5343_/A
+ sky130_fd_sc_hd__o32a_1
X_8061_ _8324_/B _8061_/B vssd1 vssd1 vccd1 vccd1 _8062_/B sky130_fd_sc_hd__nand2_2
XFILLER_126_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7012_ _7010_/X _7011_/X _7010_/X _7011_/X vssd1 vssd1 vccd1 vccd1 _7012_/X sky130_fd_sc_hd__a2bb2o_1
X_5273_ _9742_/Q _5273_/B vssd1 vssd1 vccd1 vccd1 _5273_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8963_ _8953_/X _8962_/X _8953_/X _8962_/X vssd1 vssd1 vccd1 vccd1 _8963_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8894_ _8892_/X _8893_/X _8892_/X _8893_/X vssd1 vssd1 vccd1 vccd1 _8894_/Y sky130_fd_sc_hd__o2bb2ai_1
X_7914_ _7914_/A vssd1 vssd1 vccd1 vccd1 _9507_/S sky130_fd_sc_hd__clkinv_8
XFILLER_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7845_ _9913_/Q _7841_/Y _7818_/X _7848_/B vssd1 vssd1 vccd1 vccd1 _7845_/X sky130_fd_sc_hd__o211a_1
XPHY_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4988_ _9843_/Q _4985_/X input40/X _4987_/X _4974_/X vssd1 vssd1 vccd1 vccd1 _9843_/D
+ sky130_fd_sc_hd__o221a_1
X_7776_ _7776_/A _7781_/A vssd1 vssd1 vccd1 vccd1 _7776_/Y sky130_fd_sc_hd__nor2_1
X_9515_ _9847_/Q _9028_/X _7970_/Y _9029_/X _8970_/X _9053_/S vssd1 vssd1 vccd1 vccd1
+ _9515_/X sky130_fd_sc_hd__mux4_2
XPHY_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6727_ _6716_/A _6716_/B _6716_/X vssd1 vssd1 vccd1 vccd1 _6728_/B sky130_fd_sc_hd__a21bo_1
X_9446_ _8442_/Y _8441_/B _9490_/S vssd1 vssd1 vccd1 vccd1 _9446_/X sky130_fd_sc_hd__mux2_2
XFILLER_164_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6658_ _6658_/A _6658_/B vssd1 vssd1 vccd1 vccd1 _6669_/A sky130_fd_sc_hd__or2_1
XFILLER_194_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5609_ _5609_/A _5609_/B vssd1 vssd1 vccd1 vccd1 _9704_/D sky130_fd_sc_hd__nor2_1
X_9377_ _8433_/Y _8430_/X _9477_/S vssd1 vssd1 vccd1 vccd1 _9377_/X sky130_fd_sc_hd__mux2_4
X_6589_ _6764_/A vssd1 vssd1 vccd1 vccd1 _6660_/A sky130_fd_sc_hd__clkbuf_2
X_8328_ _8328_/A _8328_/B _8328_/C _8310_/X vssd1 vssd1 vccd1 vccd1 _8331_/A sky130_fd_sc_hd__or4b_4
XFILLER_11_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8259_ _8259_/A vssd1 vssd1 vccd1 vccd1 _8259_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _9930_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput27 io_wb_dat_i[1] vssd1 vssd1 vccd1 vccd1 _5039_/A sky130_fd_sc_hd__buf_6
Xinput16 io_wb_dat_i[0] vssd1 vssd1 vccd1 vccd1 _5041_/A sky130_fd_sc_hd__buf_6
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput38 io_wb_dat_i[2] vssd1 vssd1 vccd1 vccd1 _4860_/A sky130_fd_sc_hd__buf_6
XFILLER_10_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput49 reset vssd1 vssd1 vccd1 vccd1 _5214_/A sky130_fd_sc_hd__buf_4
XFILLER_143_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5960_ _9074_/X _5958_/X _9569_/Q _5959_/X vssd1 vssd1 vccd1 vccd1 _9569_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5891_ _5891_/A vssd1 vssd1 vccd1 vccd1 _5891_/X sky130_fd_sc_hd__buf_2
X_4911_ _5586_/A vssd1 vssd1 vccd1 vccd1 _5662_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_206_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7630_ _7069_/A _7069_/B _7070_/B vssd1 vssd1 vccd1 vccd1 _7630_/Y sky130_fd_sc_hd__o21ai_1
X_4842_ _9900_/Q vssd1 vssd1 vccd1 vccd1 _7657_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4773_ _9326_/X _4763_/X _7683_/A _4767_/X _5916_/A vssd1 vssd1 vccd1 vccd1 _9926_/D
+ sky130_fd_sc_hd__o221a_1
X_7561_ _7529_/X _7554_/Y _7529_/X _7554_/Y vssd1 vssd1 vccd1 vccd1 _7578_/A sky130_fd_sc_hd__a2bb2o_1
X_6512_ _6317_/B _6409_/A _6511_/X vssd1 vssd1 vccd1 vccd1 _6512_/Y sky130_fd_sc_hd__o21ai_1
X_9300_ _9770_/Q _9299_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9300_/X sky130_fd_sc_hd__mux2_1
X_7492_ _7121_/X _7492_/B _7492_/C _7492_/D vssd1 vssd1 vccd1 vccd1 _7492_/X sky130_fd_sc_hd__and4b_2
XFILLER_173_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9231_ _7782_/Y _9750_/Q _9327_/S vssd1 vssd1 vccd1 vccd1 _9231_/X sky130_fd_sc_hd__mux2_1
X_6443_ _6443_/A vssd1 vssd1 vccd1 vccd1 _6443_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9162_ _6262_/X input31/X _9170_/S vssd1 vssd1 vccd1 vccd1 _9162_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6374_ _9756_/Q _6374_/B vssd1 vssd1 vccd1 vccd1 _6443_/A sky130_fd_sc_hd__or2_1
X_9093_ _6561_/Y _6562_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9093_/X sky130_fd_sc_hd__mux2_2
X_8113_ _8111_/Y _8112_/Y _8072_/B vssd1 vssd1 vccd1 vccd1 _8113_/Y sky130_fd_sc_hd__o21ai_1
X_5325_ _9717_/Q _9716_/Q _9718_/Q vssd1 vssd1 vccd1 vccd1 _5392_/B sky130_fd_sc_hd__and3_1
X_8044_ _8044_/A _8044_/B vssd1 vssd1 vccd1 vccd1 _8044_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5256_ _5256_/A vssd1 vssd1 vccd1 vccd1 _9747_/D sky130_fd_sc_hd__inv_2
X_5187_ _5660_/A vssd1 vssd1 vccd1 vccd1 _5187_/X sky130_fd_sc_hd__buf_2
XFILLER_68_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8946_ _8943_/X _8945_/X _8943_/X _8945_/X vssd1 vssd1 vccd1 vccd1 _8946_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_83_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8877_ _8959_/A _8958_/B _8919_/A _8955_/B vssd1 vssd1 vccd1 vccd1 _8878_/B sky130_fd_sc_hd__o22a_1
XPHY_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7828_ _4820_/X _7824_/Y _7818_/X _7831_/B vssd1 vssd1 vccd1 vccd1 _7828_/X sky130_fd_sc_hd__o211a_1
XPHY_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7759_ _7755_/X _6337_/A _4794_/X _6348_/Y _7758_/X vssd1 vssd1 vccd1 vccd1 _7772_/A
+ sky130_fd_sc_hd__o221a_1
XPHY_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9429_ _8798_/X _8796_/A _9477_/S vssd1 vssd1 vccd1 vccd1 _9429_/X sky130_fd_sc_hd__mux2_2
XFILLER_192_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5110_ _5128_/A _5108_/Y _5109_/Y _5097_/X vssd1 vssd1 vccd1 vccd1 _5111_/B sky130_fd_sc_hd__o22a_1
X_6090_ _6088_/A _6085_/X _6088_/A _6085_/X vssd1 vssd1 vccd1 vccd1 _6090_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5041_ _5041_/A vssd1 vssd1 vccd1 vccd1 _5041_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_111_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9780_ _9819_/CLK _9780_/D vssd1 vssd1 vccd1 vccd1 _9780_/Q sky130_fd_sc_hd__dfxtp_1
X_8800_ _8800_/A _8800_/B vssd1 vssd1 vccd1 vccd1 _8801_/A sky130_fd_sc_hd__or2_2
X_8731_ _8680_/X _8681_/X _8640_/Y _8682_/X vssd1 vssd1 vccd1 vccd1 _8731_/X sky130_fd_sc_hd__o22a_1
X_6992_ _6992_/A _6992_/B vssd1 vssd1 vccd1 vccd1 _6992_/X sky130_fd_sc_hd__or2_1
XFILLER_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5943_ _9156_/X _5937_/X _9580_/Q _5938_/X vssd1 vssd1 vccd1 vccd1 _9580_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8662_ _8660_/X _8661_/X _8660_/X _8661_/X vssd1 vssd1 vccd1 vccd1 _8662_/Y sky130_fd_sc_hd__a2bb2oi_2
X_5874_ _9622_/Q _5865_/A _5035_/X _5866_/A _5867_/X vssd1 vssd1 vccd1 vccd1 _9622_/D
+ sky130_fd_sc_hd__o221a_1
X_8593_ _8593_/A _8593_/B vssd1 vssd1 vccd1 vccd1 _8593_/Y sky130_fd_sc_hd__nor2_4
XFILLER_138_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4825_ _9270_/X _4822_/X _7665_/A _4824_/X _4817_/X vssd1 vssd1 vccd1 vccd1 _9908_/D
+ sky130_fd_sc_hd__o221a_1
X_7613_ _7601_/A _7601_/B _7602_/B vssd1 vssd1 vccd1 vccd1 _7613_/X sky130_fd_sc_hd__a21bo_1
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7544_ _7487_/A _7522_/B _7518_/A _7490_/B vssd1 vssd1 vccd1 vccd1 _7544_/X sky130_fd_sc_hd__o22a_1
XFILLER_193_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4756_ _4776_/A vssd1 vssd1 vccd1 vccd1 _5790_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_161_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7475_ _7438_/X _7448_/X _7438_/X _7448_/X vssd1 vssd1 vccd1 vccd1 _7475_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_161_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9214_ _9819_/Q _7645_/Y _9528_/Q vssd1 vssd1 vccd1 vccd1 _9214_/X sky130_fd_sc_hd__mux2_1
X_6426_ _9765_/Q _8223_/A _8221_/A vssd1 vssd1 vccd1 vccd1 _6427_/A sky130_fd_sc_hd__a21bo_1
XFILLER_161_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6357_ _9847_/Q vssd1 vssd1 vccd1 vccd1 _8183_/A sky130_fd_sc_hd__inv_2
X_9145_ _6157_/X _5032_/A _9148_/S vssd1 vssd1 vccd1 vccd1 _9145_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5308_ _9733_/Q _9732_/Q vssd1 vssd1 vccd1 vccd1 _5308_/Y sky130_fd_sc_hd__nor2_1
X_6288_ _6288_/A _6288_/B vssd1 vssd1 vccd1 vccd1 _6296_/A sky130_fd_sc_hd__or2_1
X_9076_ _7830_/X _9761_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9076_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8027_ _8027_/A _8033_/B vssd1 vssd1 vccd1 vccd1 _8027_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5239_ _9735_/Q vssd1 vssd1 vccd1 vccd1 _5240_/C sky130_fd_sc_hd__inv_2
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8929_ _8926_/X _8928_/Y _8926_/X _8928_/Y vssd1 vssd1 vccd1 vccd1 _8930_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_140_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5590_ _5586_/X _5587_/Y _5588_/X _7646_/A _5577_/X vssd1 vssd1 vccd1 vccd1 _5591_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7260_ _7260_/A _7260_/B vssd1 vssd1 vccd1 vccd1 _7427_/B sky130_fd_sc_hd__nor2_2
XFILLER_171_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7191_ _7191_/A _7191_/B vssd1 vssd1 vccd1 vccd1 _7502_/B sky130_fd_sc_hd__nor2_2
X_6211_ _9577_/Q _6167_/A _8005_/A _6201_/A vssd1 vssd1 vccd1 vccd1 _6221_/C sky130_fd_sc_hd__a22o_1
X_6142_ _6142_/A vssd1 vssd1 vccd1 vccd1 _6193_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6073_ _9646_/Q vssd1 vssd1 vccd1 vccd1 _6074_/B sky130_fd_sc_hd__inv_2
X_9901_ _9917_/CLK _9901_/D vssd1 vssd1 vccd1 vccd1 _9901_/Q sky130_fd_sc_hd__dfxtp_2
X_5024_ _5036_/A vssd1 vssd1 vccd1 vccd1 _5024_/X sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_18 _5029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9832_ _9833_/CLK _9832_/D vssd1 vssd1 vccd1 vccd1 _9832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6975_ _6975_/A _9465_/X vssd1 vssd1 vccd1 vccd1 _6975_/X sky130_fd_sc_hd__or2_1
X_9763_ _9915_/CLK _9763_/D vssd1 vssd1 vccd1 vccd1 _9763_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5926_ _9169_/X _5921_/X _9593_/Q _5924_/X vssd1 vssd1 vccd1 vccd1 _9593_/D sky130_fd_sc_hd__a22o_1
XFILLER_179_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8714_ _8714_/A vssd1 vssd1 vccd1 vccd1 _8714_/Y sky130_fd_sc_hd__inv_2
X_9694_ _9699_/CLK _9694_/D vssd1 vssd1 vccd1 vccd1 _9694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8645_ _8645_/A _8645_/B vssd1 vssd1 vccd1 vccd1 _8695_/A sky130_fd_sc_hd__or2_1
XFILLER_110_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5857_ _9629_/Q _5847_/A _4860_/X _5848_/A _5853_/X vssd1 vssd1 vccd1 vccd1 _9629_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_139_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8576_ _8576_/A _8766_/B _8576_/C vssd1 vssd1 vccd1 vccd1 _8576_/X sky130_fd_sc_hd__or3_1
XFILLER_194_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4808_ _9083_/X _4796_/X _9914_/Q _4799_/X _4806_/X vssd1 vssd1 vccd1 vccd1 _9914_/D
+ sky130_fd_sc_hd__o221a_1
X_5788_ _6558_/A _9658_/Q _5731_/Y vssd1 vssd1 vccd1 vccd1 _5788_/X sky130_fd_sc_hd__a21o_1
XFILLER_135_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7527_ _7263_/X _7482_/X _7263_/X _7482_/X vssd1 vssd1 vccd1 vccd1 _7527_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7458_ _7457_/A _7457_/B _7457_/X vssd1 vssd1 vccd1 vccd1 _7470_/A sky130_fd_sc_hd__a21boi_2
X_6409_ _6409_/A vssd1 vssd1 vccd1 vccd1 _6545_/B sky130_fd_sc_hd__inv_2
XFILLER_134_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7389_ _7389_/A _7389_/B vssd1 vssd1 vccd1 vccd1 _7467_/A sky130_fd_sc_hd__or2_1
XFILLER_115_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9128_ _9865_/Q _9881_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9128_/X sky130_fd_sc_hd__mux2_1
X_9059_ _8026_/Y _8024_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9059_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6760_ _6760_/A _6760_/B _6760_/C vssd1 vssd1 vccd1 vccd1 _6760_/X sky130_fd_sc_hd__or3_4
XFILLER_35_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5711_ _5041_/A _5710_/A _9667_/Q _5710_/Y _5698_/X vssd1 vssd1 vccd1 vccd1 _9667_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_62_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6691_ _6713_/A _6691_/B _6691_/C vssd1 vssd1 vccd1 vccd1 _6995_/A sky130_fd_sc_hd__and3_1
XFILLER_148_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8430_ _8432_/A _8398_/X _8432_/A _8398_/X vssd1 vssd1 vccd1 vccd1 _8430_/X sky130_fd_sc_hd__a2bb2o_1
X_5642_ _9679_/Q vssd1 vssd1 vccd1 vccd1 _6578_/A sky130_fd_sc_hd__clkbuf_2
X_8361_ _4780_/X _8359_/Y _7682_/A _8354_/Y _8360_/X vssd1 vssd1 vccd1 vccd1 _8361_/X
+ sky130_fd_sc_hd__o221a_1
X_5573_ _5573_/A vssd1 vssd1 vccd1 vccd1 _5573_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7312_ _7312_/A _7311_/X vssd1 vssd1 vccd1 vccd1 _7312_/X sky130_fd_sc_hd__or2b_1
X_8292_ _7877_/A _8210_/X _7882_/A _8208_/Y _8291_/X vssd1 vssd1 vccd1 vccd1 _8292_/X
+ sky130_fd_sc_hd__o221a_1
X_7243_ _7243_/A _7222_/X vssd1 vssd1 vccd1 vccd1 _7245_/A sky130_fd_sc_hd__or2b_1
X_7174_ _7174_/A _7153_/X vssd1 vssd1 vccd1 vccd1 _7176_/A sky130_fd_sc_hd__or2b_1
XFILLER_112_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6125_ _9565_/Q vssd1 vssd1 vccd1 vccd1 _6125_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6056_ _6056_/A _6056_/B vssd1 vssd1 vccd1 vccd1 _6057_/A sky130_fd_sc_hd__or2_2
XFILLER_85_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5007_ _9831_/Q _5003_/X input26/X _5004_/X _5000_/X vssd1 vssd1 vccd1 vccd1 _9831_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9815_ _9819_/CLK _9815_/D vssd1 vssd1 vccd1 vccd1 _9815_/Q sky130_fd_sc_hd__dfxtp_1
X_9746_ _9893_/CLK _9746_/D vssd1 vssd1 vccd1 vccd1 _9746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6958_ _6933_/X _6937_/X _6938_/X _6957_/Y vssd1 vssd1 vccd1 vccd1 _6958_/X sky130_fd_sc_hd__o22a_1
XFILLER_53_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9677_ _9699_/CLK _9677_/D vssd1 vssd1 vccd1 vccd1 _9677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5909_ _5909_/A _9133_/X vssd1 vssd1 vccd1 vccd1 _9601_/D sky130_fd_sc_hd__and2_1
X_6889_ _6876_/X _6877_/X _6876_/X _6877_/X vssd1 vssd1 vccd1 vccd1 _6889_/X sky130_fd_sc_hd__a2bb2o_2
X_8628_ _8628_/A _8586_/X vssd1 vssd1 vccd1 vccd1 _8629_/A sky130_fd_sc_hd__or2b_1
XFILLER_167_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8559_ _8559_/A _8559_/B vssd1 vssd1 vccd1 vccd1 _8603_/A sky130_fd_sc_hd__nand2_1
XFILLER_139_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7930_ _9485_/X _7956_/B vssd1 vssd1 vccd1 vccd1 _7930_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7861_ _7861_/A _7861_/B vssd1 vssd1 vccd1 vccd1 _7865_/B sky130_fd_sc_hd__or2_2
XFILLER_63_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6812_ _6812_/A _6862_/A vssd1 vssd1 vccd1 vccd1 _6813_/A sky130_fd_sc_hd__or2_2
X_9600_ _9895_/CLK _9600_/D vssd1 vssd1 vccd1 vccd1 _9600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7792_ _7793_/A _7658_/B _7659_/B vssd1 vssd1 vccd1 vccd1 _7792_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_63_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9531_ _9796_/CLK _9531_/D vssd1 vssd1 vccd1 vccd1 _9531_/Q sky130_fd_sc_hd__dfxtp_1
X_6743_ _6743_/A _6743_/B vssd1 vssd1 vccd1 vccd1 _6910_/B sky130_fd_sc_hd__nor2_2
X_9462_ _5721_/X _6581_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9462_/X sky130_fd_sc_hd__mux2_2
X_6674_ _6674_/A _6991_/B vssd1 vssd1 vccd1 vccd1 _6674_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5625_ _8176_/A _5625_/B vssd1 vssd1 vccd1 vccd1 _9701_/D sky130_fd_sc_hd__nor2_1
XFILLER_149_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8413_ _9699_/Q _9683_/Q _8412_/Y _6982_/C vssd1 vssd1 vccd1 vccd1 _8413_/X sky130_fd_sc_hd__o22a_2
XFILLER_164_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9393_ _8744_/X _8742_/A _9490_/S vssd1 vssd1 vccd1 vccd1 _9393_/X sky130_fd_sc_hd__mux2_2
X_8344_ _7673_/A _8342_/Y _4802_/X _8337_/Y _8343_/X vssd1 vssd1 vccd1 vccd1 _8344_/X
+ sky130_fd_sc_hd__o221a_1
X_5556_ _9714_/Q vssd1 vssd1 vccd1 vccd1 _7652_/A sky130_fd_sc_hd__inv_2
XFILLER_117_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8275_ _9910_/Q _8233_/Y _8274_/Y vssd1 vssd1 vccd1 vccd1 _8275_/X sky130_fd_sc_hd__o21ba_1
XFILLER_2_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5487_ _5419_/X _5458_/X _5419_/X _5458_/X vssd1 vssd1 vccd1 vccd1 _5487_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7226_ _7385_/A _7238_/B vssd1 vssd1 vccd1 vccd1 _7234_/C sky130_fd_sc_hd__nor2_1
XFILLER_120_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7157_ _7155_/X _7156_/X _7155_/X _7156_/X vssd1 vssd1 vccd1 vccd1 _7164_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_112_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6108_ _9862_/Q _6101_/Y _6103_/A _6105_/X vssd1 vssd1 vccd1 vccd1 _6108_/X sky130_fd_sc_hd__o22a_1
XFILLER_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7088_ _7088_/A _7088_/B vssd1 vssd1 vccd1 vccd1 _7089_/B sky130_fd_sc_hd__or2_1
X_6039_ _7962_/A _9641_/Q _6026_/Y _6031_/A vssd1 vssd1 vccd1 vccd1 _6039_/X sky130_fd_sc_hd__o22a_1
XFILLER_100_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9729_ _9874_/CLK _9729_/D vssd1 vssd1 vccd1 vccd1 _9729_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6390_ _9772_/Q _6390_/B vssd1 vssd1 vccd1 vccd1 _8203_/A sky130_fd_sc_hd__or2_2
X_5410_ _9348_/X vssd1 vssd1 vccd1 vccd1 _5412_/A sky130_fd_sc_hd__inv_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5341_ _9335_/X _5692_/A _5340_/X vssd1 vssd1 vccd1 vccd1 _5341_/Y sky130_fd_sc_hd__a21oi_1
X_8060_ _4960_/X _8050_/Y _8051_/Y _8059_/X vssd1 vssd1 vccd1 vccd1 _8061_/B sky130_fd_sc_hd__o22a_1
XFILLER_141_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7011_ _6998_/X _7003_/X _6998_/X _7003_/X vssd1 vssd1 vccd1 vccd1 _7011_/X sky130_fd_sc_hd__a2bb2o_1
X_5272_ _5272_/A vssd1 vssd1 vccd1 vccd1 _5273_/B sky130_fd_sc_hd__inv_2
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8962_ _8956_/X _8961_/Y _8956_/X _8961_/Y vssd1 vssd1 vccd1 vccd1 _8962_/X sky130_fd_sc_hd__a2bb2o_1
X_7913_ _7913_/A vssd1 vssd1 vccd1 vccd1 _9506_/S sky130_fd_sc_hd__clkinv_8
XFILLER_55_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8893_ _8955_/A _8893_/B _8893_/C vssd1 vssd1 vccd1 vccd1 _8893_/X sky130_fd_sc_hd__or3_4
X_7844_ _7844_/A _7844_/B vssd1 vssd1 vccd1 vccd1 _7848_/B sky130_fd_sc_hd__or2_2
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7775_ _7839_/A vssd1 vssd1 vccd1 vccd1 _7781_/A sky130_fd_sc_hd__buf_4
XPHY_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4987_ _5004_/A vssd1 vssd1 vccd1 vccd1 _4987_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6726_ _6726_/A _6705_/X vssd1 vssd1 vccd1 vccd1 _6728_/A sky130_fd_sc_hd__or2b_1
X_9514_ _9846_/Q _9025_/X _7964_/Y _9026_/X _8970_/X _9053_/S vssd1 vssd1 vccd1 vccd1
+ _9514_/X sky130_fd_sc_hd__mux4_2
XPHY_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6657_ _6646_/A _6646_/B _6646_/X vssd1 vssd1 vccd1 vccd1 _6658_/B sky130_fd_sc_hd__a21bo_1
X_9445_ _9526_/Q _5039_/A _9445_/S vssd1 vssd1 vccd1 vccd1 _9445_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5608_ _5586_/X _5604_/Y _5605_/Y _7640_/A _5607_/X vssd1 vssd1 vccd1 vccd1 _5609_/B
+ sky130_fd_sc_hd__o32a_1
X_9376_ _9291_/S _7773_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9376_/X sky130_fd_sc_hd__mux2_1
X_6588_ _6812_/A vssd1 vssd1 vccd1 vccd1 _6764_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_191_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8327_ _8369_/C _8325_/Y _8369_/B vssd1 vssd1 vccd1 vccd1 _8327_/X sky130_fd_sc_hd__a21bo_1
X_5539_ _9393_/X _5485_/X _5573_/A vssd1 vssd1 vccd1 vccd1 _5539_/X sky130_fd_sc_hd__o21a_1
XFILLER_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8258_ _8252_/X _8257_/X _8134_/A _8257_/B vssd1 vssd1 vccd1 vccd1 _8259_/A sky130_fd_sc_hd__a22o_1
XFILLER_160_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8189_ _9846_/Q _6364_/Y _8184_/Y _8188_/Y vssd1 vssd1 vccd1 vccd1 _8189_/X sky130_fd_sc_hd__o22a_1
XFILLER_160_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7209_ _7148_/X _7208_/X _7148_/X _7208_/X vssd1 vssd1 vccd1 vccd1 _7209_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_59_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput28 io_wb_dat_i[20] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput17 io_wb_dat_i[10] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_4
XFILLER_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput39 io_wb_dat_i[30] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_4
XPHY_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5890_ _9615_/Q vssd1 vssd1 vccd1 vccd1 _5890_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4910_ _9873_/Q _4905_/X _9725_/Q _4903_/X _4906_/X vssd1 vssd1 vccd1 vccd1 _9873_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4841_ _9242_/X _4834_/X _8324_/A _4836_/X _4830_/X vssd1 vssd1 vccd1 vccd1 _9901_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4772_ _9926_/Q vssd1 vssd1 vccd1 vccd1 _7683_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_193_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7560_ _7560_/A vssd1 vssd1 vccd1 vccd1 _7560_/X sky130_fd_sc_hd__buf_1
XFILLER_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6511_ _6317_/C _6411_/Y _6510_/X vssd1 vssd1 vccd1 vccd1 _6511_/X sky130_fd_sc_hd__a21o_1
XFILLER_158_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7491_ _7491_/A _7491_/B vssd1 vssd1 vccd1 vccd1 _7491_/X sky130_fd_sc_hd__or2_1
X_9230_ _9229_/X _5039_/A _9334_/S vssd1 vssd1 vccd1 vccd1 _9230_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6442_ _9791_/Q _6527_/B vssd1 vssd1 vccd1 vccd1 _6463_/B sky130_fd_sc_hd__nor2_1
XFILLER_161_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9161_ _6258_/Y input30/X _9170_/S vssd1 vssd1 vccd1 vccd1 _9161_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6373_ _9755_/Q _6467_/A vssd1 vssd1 vccd1 vccd1 _6374_/B sky130_fd_sc_hd__or2_2
XFILLER_114_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8112_ _8112_/A vssd1 vssd1 vccd1 vccd1 _8112_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9092_ _6551_/Y _6560_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9092_/X sky130_fd_sc_hd__mux2_1
X_5324_ _9720_/Q vssd1 vssd1 vccd1 vccd1 _5327_/A sky130_fd_sc_hd__inv_2
X_8043_ _8994_/X _8045_/B vssd1 vssd1 vccd1 vccd1 _8043_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5255_ _9747_/Q _5224_/X _5251_/Y _5252_/Y _5258_/A vssd1 vssd1 vccd1 vccd1 _5256_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_102_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5186_ _9764_/Q vssd1 vssd1 vccd1 vccd1 _6353_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8945_ _8862_/X _8944_/Y _8862_/X _8944_/Y vssd1 vssd1 vccd1 vccd1 _8945_/X sky130_fd_sc_hd__a2bb2o_1
X_8876_ _8876_/A vssd1 vssd1 vccd1 vccd1 _8878_/A sky130_fd_sc_hd__inv_2
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7827_ _7827_/A _7827_/B vssd1 vssd1 vccd1 vccd1 _7831_/B sky130_fd_sc_hd__or2_2
XFILLER_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7758_ _7906_/A _9778_/Q _8174_/A _9779_/Q vssd1 vssd1 vccd1 vccd1 _7758_/X sky130_fd_sc_hd__o22a_2
XPHY_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7689_ _4847_/X _6364_/Y _7793_/A _9752_/Q vssd1 vssd1 vccd1 vccd1 _7689_/X sky130_fd_sc_hd__o22a_1
X_6709_ _6868_/A _6721_/B vssd1 vssd1 vccd1 vccd1 _6717_/C sky130_fd_sc_hd__nor2_1
XPHY_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9428_ _8600_/X _8598_/Y _9490_/S vssd1 vssd1 vccd1 vccd1 _9428_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9359_ _7619_/X _7584_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9359_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5040_ _9813_/Q _5003_/A _5039_/X _5004_/A _5036_/X vssd1 vssd1 vccd1 vccd1 _9813_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_97_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6991_ _6991_/A _6991_/B vssd1 vssd1 vccd1 vccd1 _6992_/B sky130_fd_sc_hd__nor2_1
X_8730_ _8728_/X _8729_/X _8728_/X _8729_/X vssd1 vssd1 vccd1 vccd1 _8730_/X sky130_fd_sc_hd__a2bb2o_1
X_5942_ _9157_/X _5937_/X _9581_/Q _5938_/X vssd1 vssd1 vccd1 vccd1 _9581_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8661_ _8535_/X _8614_/A _8735_/A _8768_/A vssd1 vssd1 vccd1 vccd1 _8661_/X sky130_fd_sc_hd__a211o_1
X_5873_ _5872_/X _5865_/X _4978_/A _5866_/X _5867_/X vssd1 vssd1 vccd1 vccd1 _9623_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8592_ _8591_/A _8591_/B _8715_/A vssd1 vssd1 vccd1 vccd1 _8593_/B sky130_fd_sc_hd__a21o_1
X_4824_ _4836_/A vssd1 vssd1 vccd1 vccd1 _4824_/X sky130_fd_sc_hd__clkbuf_2
X_7612_ _7078_/A _7078_/B _7079_/B vssd1 vssd1 vccd1 vccd1 _7612_/X sky130_fd_sc_hd__a21bo_1
XFILLER_33_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4755_ _5214_/A vssd1 vssd1 vccd1 vccd1 _4776_/A sky130_fd_sc_hd__inv_2
XFILLER_21_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7543_ _7454_/X _7473_/Y _7454_/X _7473_/Y vssd1 vssd1 vccd1 vccd1 _7543_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_193_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9213_ _9818_/Q _7643_/Y _9528_/Q vssd1 vssd1 vccd1 vccd1 _9213_/X sky130_fd_sc_hd__mux2_1
X_7474_ _7449_/X _7453_/X _7454_/X _7473_/Y vssd1 vssd1 vccd1 vccd1 _7474_/X sky130_fd_sc_hd__o22a_1
X_6425_ _6351_/A _8221_/A _8219_/A vssd1 vssd1 vccd1 vccd1 _6428_/A sky130_fd_sc_hd__a21bo_1
XFILLER_119_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6356_ _9752_/Q vssd1 vssd1 vccd1 vccd1 _8191_/A sky130_fd_sc_hd__inv_2
XFILLER_108_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9144_ _6153_/Y _4978_/A _9148_/S vssd1 vssd1 vccd1 vccd1 _9144_/X sky130_fd_sc_hd__mux2_1
X_9075_ _6131_/X _4860_/A _9155_/S vssd1 vssd1 vccd1 vccd1 _9075_/X sky130_fd_sc_hd__mux2_1
X_5307_ _4853_/X _5240_/A _5306_/X vssd1 vssd1 vccd1 vccd1 _9734_/D sky130_fd_sc_hd__o21ai_1
X_6287_ _6268_/X _6271_/X _6285_/X _6276_/X _6286_/X vssd1 vssd1 vccd1 vccd1 _6288_/B
+ sky130_fd_sc_hd__o311a_1
X_8026_ _9071_/X _8037_/B vssd1 vssd1 vccd1 vccd1 _8026_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5238_ _5238_/A _5238_/B vssd1 vssd1 vccd1 vccd1 _5305_/A sky130_fd_sc_hd__or2_2
X_5169_ _9773_/Q _5167_/X input33/X _5168_/X _5165_/X vssd1 vssd1 vccd1 vccd1 _9773_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_124_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8928_ _8847_/Y _8927_/Y _8883_/Y vssd1 vssd1 vccd1 vccd1 _8928_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8859_ _8859_/A _8859_/B vssd1 vssd1 vccd1 vccd1 _8859_/X sky130_fd_sc_hd__or2_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7190_ _7190_/A _7190_/B vssd1 vssd1 vccd1 vccd1 _7191_/B sky130_fd_sc_hd__or2_2
X_6210_ _9577_/Q vssd1 vssd1 vccd1 vccd1 _8005_/A sky130_fd_sc_hd__inv_2
X_6141_ _6141_/A vssd1 vssd1 vccd1 vccd1 _6142_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6072_ _6066_/Y _6071_/A _6066_/A _6071_/Y vssd1 vssd1 vccd1 vccd1 _6072_/X sky130_fd_sc_hd__o22a_1
X_9900_ _9903_/CLK _9900_/D vssd1 vssd1 vccd1 vccd1 _9900_/Q sky130_fd_sc_hd__dfxtp_1
X_5023_ _9821_/Q _5019_/X input47/X _5020_/X _5016_/X vssd1 vssd1 vccd1 vccd1 _9821_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_38_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_19 _5026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_9831_ _9833_/CLK _9831_/D vssd1 vssd1 vccd1 vccd1 _9831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6974_ _6978_/C _9467_/X vssd1 vssd1 vccd1 vccd1 _6974_/Y sky130_fd_sc_hd__nor2_1
X_9762_ _9915_/CLK _9762_/D vssd1 vssd1 vccd1 vccd1 _9762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5925_ _9170_/X _5921_/X _9594_/Q _5924_/X vssd1 vssd1 vccd1 vccd1 _9594_/D sky130_fd_sc_hd__a22o_1
XFILLER_179_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8713_ _8711_/X _8712_/X _8711_/X _8712_/X vssd1 vssd1 vccd1 vccd1 _8713_/X sky130_fd_sc_hd__a2bb2o_1
X_9693_ _9699_/CLK _9693_/D vssd1 vssd1 vccd1 vccd1 _9693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5856_ _8823_/A _5847_/X _5035_/X _5848_/X _5853_/X vssd1 vssd1 vccd1 vccd1 _9630_/D
+ sky130_fd_sc_hd__o221a_1
X_8644_ _8644_/A vssd1 vssd1 vccd1 vccd1 _8645_/B sky130_fd_sc_hd__inv_2
XFILLER_139_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4807_ _9290_/X _4796_/X _9915_/Q _4799_/X _4806_/X vssd1 vssd1 vccd1 vccd1 _9915_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8575_ _8584_/B vssd1 vssd1 vccd1 vccd1 _8766_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_166_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5787_ _5787_/A vssd1 vssd1 vccd1 vccd1 _5787_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7526_ _7489_/X _7525_/Y _7489_/X _7525_/Y vssd1 vssd1 vccd1 vccd1 _7526_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_147_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7457_ _7457_/A _7457_/B vssd1 vssd1 vccd1 vccd1 _7457_/X sky130_fd_sc_hd__or2_2
X_6408_ _6345_/Y _6407_/Y _6393_/B vssd1 vssd1 vccd1 vccd1 _6409_/A sky130_fd_sc_hd__o21ai_2
XFILLER_162_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9127_ _9864_/Q _9880_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9127_/X sky130_fd_sc_hd__mux2_1
X_7388_ _7389_/A _7398_/B vssd1 vssd1 vccd1 vccd1 _7394_/C sky130_fd_sc_hd__nor2_1
X_6339_ _9757_/Q vssd1 vssd1 vccd1 vccd1 _6339_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9058_ _8022_/Y _8021_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9058_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8009_ _9413_/X _8009_/B vssd1 vssd1 vccd1 vccd1 _8009_/Y sky130_fd_sc_hd__nor2_1
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5710_ _5710_/A vssd1 vssd1 vccd1 vccd1 _5710_/Y sky130_fd_sc_hd__inv_2
X_6690_ _6623_/X _6689_/X _6623_/X _6689_/X vssd1 vssd1 vccd1 vccd1 _6690_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5641_ _9696_/Q _5631_/X _6596_/A _5635_/X _5632_/X vssd1 vssd1 vccd1 vccd1 _9696_/D
+ sky130_fd_sc_hd__o221a_1
X_8360_ _7892_/A _9556_/Q _7885_/X _9555_/Q vssd1 vssd1 vccd1 vccd1 _8360_/X sky130_fd_sc_hd__o22a_1
X_5572_ _9711_/Q _4922_/X _5570_/X _5571_/Y _5187_/X vssd1 vssd1 vccd1 vccd1 _9711_/D
+ sky130_fd_sc_hd__o221a_1
X_8291_ _7877_/A _8210_/X _7728_/X _8212_/Y _8290_/X vssd1 vssd1 vccd1 vccd1 _8291_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_117_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7311_ _7311_/A _7385_/B _7331_/A _7379_/A vssd1 vssd1 vccd1 vccd1 _7311_/X sky130_fd_sc_hd__or4_4
XFILLER_144_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7242_ _7247_/A _7222_/B _7400_/A _7247_/B vssd1 vssd1 vccd1 vccd1 _7243_/A sky130_fd_sc_hd__o22a_1
XFILLER_116_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7173_ _7290_/A _9430_/X _7265_/A _7178_/B vssd1 vssd1 vccd1 vccd1 _7174_/A sky130_fd_sc_hd__o22a_1
XFILLER_131_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6124_ _9563_/Q _6123_/X _9563_/Q _6123_/X vssd1 vssd1 vccd1 vccd1 _6124_/X sky130_fd_sc_hd__o2bb2a_1
X_6055_ _9857_/Q _6055_/B vssd1 vssd1 vccd1 vccd1 _6056_/B sky130_fd_sc_hd__nor2_1
X_5006_ _9832_/Q _5003_/X input28/X _5004_/X _5000_/X vssd1 vssd1 vccd1 vccd1 _9832_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_66_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9814_ _9819_/CLK _9814_/D vssd1 vssd1 vccd1 vccd1 _9814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9745_ _9887_/CLK _9745_/D vssd1 vssd1 vccd1 vccd1 _9745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6957_ _6957_/A vssd1 vssd1 vccd1 vccd1 _6957_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9676_ _9699_/CLK _9676_/D vssd1 vssd1 vccd1 vccd1 _9676_/Q sky130_fd_sc_hd__dfxtp_2
X_5908_ _5909_/A _9134_/X vssd1 vssd1 vccd1 vccd1 _9602_/D sky130_fd_sc_hd__and2_1
X_6888_ _6888_/A _6888_/B vssd1 vssd1 vccd1 vccd1 _6899_/A sky130_fd_sc_hd__or2_1
XFILLER_194_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8627_ _8766_/C _8626_/X _8766_/C _8626_/X vssd1 vssd1 vccd1 vccd1 _8627_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_179_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5839_ _4860_/X _5818_/X _9637_/Q _5819_/X _5070_/A vssd1 vssd1 vccd1 vccd1 _9637_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8558_ _8403_/X _8557_/X _8403_/X _8557_/X vssd1 vssd1 vccd1 vccd1 _8559_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_182_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7509_ _7498_/X _7508_/X _7498_/X _7508_/X vssd1 vssd1 vccd1 vccd1 _7509_/X sky130_fd_sc_hd__a2bb2o_1
X_8489_ _8401_/Y _8488_/X _8401_/Y _8488_/X vssd1 vssd1 vccd1 vccd1 _8491_/B sky130_fd_sc_hd__a2bb2o_2
XFILLER_107_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7860_ _7860_/A vssd1 vssd1 vccd1 vccd1 _7860_/X sky130_fd_sc_hd__buf_2
X_6811_ _6868_/B vssd1 vssd1 vccd1 vccd1 _6883_/B sky130_fd_sc_hd__buf_1
X_7791_ _7788_/A _7788_/B _7789_/Y _7790_/X vssd1 vssd1 vccd1 vccd1 _7791_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_196_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9530_ _9898_/CLK _9530_/D vssd1 vssd1 vccd1 vccd1 _9530_/Q sky130_fd_sc_hd__dfxtp_2
X_6742_ _6742_/A _6742_/B vssd1 vssd1 vccd1 vccd1 _6743_/B sky130_fd_sc_hd__or2_2
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9461_ _5717_/Y _6580_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9461_/X sky130_fd_sc_hd__mux2_1
X_6673_ _6673_/A _6673_/B vssd1 vssd1 vccd1 vccd1 _6991_/B sky130_fd_sc_hd__nor2_2
XFILLER_176_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5624_ _5704_/A _5621_/Y _5622_/X _7637_/A _5607_/X vssd1 vssd1 vccd1 vccd1 _5625_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_149_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9392_ _8604_/X _8602_/A _9477_/S vssd1 vssd1 vccd1 vccd1 _9392_/X sky130_fd_sc_hd__mux2_1
X_8412_ _9699_/Q vssd1 vssd1 vccd1 vccd1 _8412_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8343_ _7692_/X _9548_/Q _7738_/X _9547_/Q vssd1 vssd1 vccd1 vccd1 _8343_/X sky130_fd_sc_hd__o22a_1
X_5555_ _5555_/A _5555_/B vssd1 vssd1 vccd1 vccd1 _5555_/Y sky130_fd_sc_hd__nor2_1
XFILLER_172_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5486_ _9393_/X _5485_/X _9393_/X _5485_/X vssd1 vssd1 vccd1 vccd1 _5574_/A sky130_fd_sc_hd__a2bb2oi_1
X_8274_ _7666_/A _8234_/Y _8273_/Y vssd1 vssd1 vccd1 vccd1 _8274_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7225_ _7223_/X _7224_/X _7223_/X _7224_/X vssd1 vssd1 vccd1 vccd1 _7233_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_132_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7156_ _7156_/A _9424_/X vssd1 vssd1 vccd1 vccd1 _7156_/X sky130_fd_sc_hd__or2_1
XFILLER_112_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6107_ _6103_/X _6104_/X _6103_/X _6104_/X vssd1 vssd1 vccd1 vccd1 _6107_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7087_ _7087_/A _7087_/B vssd1 vssd1 vccd1 vccd1 _7088_/B sky130_fd_sc_hd__or2_1
XFILLER_58_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6038_ _6036_/Y _6037_/X _6036_/Y _6037_/X vssd1 vssd1 vccd1 vccd1 _6038_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7989_ _8986_/X _8002_/B vssd1 vssd1 vccd1 vccd1 _7989_/Y sky130_fd_sc_hd__nor2_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9728_ _9874_/CLK _9728_/D vssd1 vssd1 vccd1 vccd1 _9728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9659_ _9673_/CLK _9659_/D vssd1 vssd1 vccd1 vccd1 _9659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5340_ _5919_/A _5586_/A _5340_/C vssd1 vssd1 vccd1 vccd1 _5340_/X sky130_fd_sc_hd__and3_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5271_ _5271_/A vssd1 vssd1 vccd1 vccd1 _5271_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_141_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7010_ _6746_/X _6964_/X _6746_/X _6964_/X vssd1 vssd1 vccd1 vccd1 _7010_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_141_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8961_ _8957_/Y _8960_/X _8957_/Y _8960_/X vssd1 vssd1 vccd1 vccd1 _8961_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7912_ _7912_/A vssd1 vssd1 vccd1 vccd1 _9505_/S sky130_fd_sc_hd__clkinv_8
XFILLER_95_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8892_ _8774_/A _8851_/A _8852_/X _8853_/X vssd1 vssd1 vccd1 vccd1 _8892_/X sky130_fd_sc_hd__o22a_1
XFILLER_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7843_ _7743_/X _7837_/Y _7671_/B vssd1 vssd1 vccd1 vccd1 _7843_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_36_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4986_ _5030_/A vssd1 vssd1 vccd1 vccd1 _5004_/A sky130_fd_sc_hd__clkbuf_4
X_7774_ _7773_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _7839_/A sky130_fd_sc_hd__nand2b_4
XPHY_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6725_ _6730_/A _6705_/B _6883_/A _6730_/B vssd1 vssd1 vccd1 vccd1 _6726_/A sky130_fd_sc_hd__o22a_1
X_9513_ _9845_/Q _9022_/X _7956_/Y _9023_/X _8970_/X _9053_/S vssd1 vssd1 vccd1 vccd1
+ _9513_/X sky130_fd_sc_hd__mux4_2
XPHY_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6656_ _6656_/A _6632_/X vssd1 vssd1 vccd1 vccd1 _6658_/A sky130_fd_sc_hd__or2b_1
X_9444_ _9527_/Q _4860_/A _9445_/S vssd1 vssd1 vccd1 vccd1 _9444_/X sky130_fd_sc_hd__mux2_1
X_5607_ _5644_/A vssd1 vssd1 vccd1 vccd1 _5607_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_9375_ _9374_/X _7005_/A _9507_/S vssd1 vssd1 vccd1 vccd1 _9375_/X sky130_fd_sc_hd__mux2_1
X_6587_ _6821_/B vssd1 vssd1 vccd1 vccd1 _6812_/A sky130_fd_sc_hd__buf_1
X_8326_ _7803_/A _9535_/Q _7797_/A _9534_/Q vssd1 vssd1 vccd1 vccd1 _8369_/B sky130_fd_sc_hd__a22oi_1
X_5538_ _5574_/A _5574_/B vssd1 vssd1 vccd1 vccd1 _5573_/A sky130_fd_sc_hd__nand2_1
XFILLER_191_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8257_ _8257_/A _8257_/B vssd1 vssd1 vccd1 vccd1 _8257_/X sky130_fd_sc_hd__or2_1
XFILLER_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5469_ _5406_/X _5463_/X _5406_/X _5463_/X vssd1 vssd1 vccd1 vccd1 _5469_/X sky130_fd_sc_hd__a2bb2o_2
X_7208_ _7194_/X _7205_/X _7206_/X _7207_/X vssd1 vssd1 vccd1 vccd1 _7208_/X sky130_fd_sc_hd__o22a_1
X_8188_ _6365_/Y _5218_/X _8187_/Y vssd1 vssd1 vccd1 vccd1 _8188_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_120_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7139_ _9625_/Q _7135_/Y _5872_/X _7137_/Y _7138_/X vssd1 vssd1 vccd1 vccd1 _7147_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_59_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 io_wb_dat_i[11] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_4
XFILLER_168_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput29 io_wb_dat_i[21] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_4
XFILLER_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4840_ _9901_/Q vssd1 vssd1 vccd1 vccd1 _8324_/A sky130_fd_sc_hd__clkbuf_2
X_4771_ _9330_/X _4763_/X _4770_/X _4767_/X _5916_/A vssd1 vssd1 vccd1 vccd1 _9927_/D
+ sky130_fd_sc_hd__o221a_1
X_6510_ _6317_/C _6411_/Y _6317_/D _6416_/A _6509_/Y vssd1 vssd1 vccd1 vccd1 _6510_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7490_ _7490_/A _7490_/B vssd1 vssd1 vccd1 vccd1 _7490_/X sky130_fd_sc_hd__or2_1
XFILLER_158_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6441_ _5198_/X _6377_/B _8231_/A vssd1 vssd1 vccd1 vccd1 _6527_/B sky130_fd_sc_hd__a21boi_2
X_9160_ _6253_/X input29/X _9170_/S vssd1 vssd1 vccd1 vccd1 _9160_/X sky130_fd_sc_hd__mux2_1
X_6372_ _9754_/Q _6372_/B vssd1 vssd1 vccd1 vccd1 _6467_/A sky130_fd_sc_hd__or2_1
XFILLER_161_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8111_ _9543_/Q vssd1 vssd1 vccd1 vccd1 _8111_/Y sky130_fd_sc_hd__inv_2
X_5323_ _9721_/Q vssd1 vssd1 vccd1 vccd1 _5328_/A sky130_fd_sc_hd__inv_2
X_9091_ _9090_/X input26/X _9294_/S vssd1 vssd1 vccd1 vccd1 _9091_/X sky130_fd_sc_hd__mux2_1
X_8042_ _8042_/A _8044_/B vssd1 vssd1 vccd1 vccd1 _8042_/Y sky130_fd_sc_hd__nor2_1
X_5254_ _5251_/Y _5253_/Y _5222_/A vssd1 vssd1 vccd1 vccd1 _5258_/A sky130_fd_sc_hd__a21oi_1
X_5185_ _9765_/Q _5178_/X input24/X _5179_/X _5175_/X vssd1 vssd1 vccd1 vccd1 _9765_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_56_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8944_ _8944_/A _8944_/B _8944_/C _9477_/S vssd1 vssd1 vccd1 vccd1 _8944_/Y sky130_fd_sc_hd__nor4_2
XFILLER_113_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8875_ _8875_/A _8958_/B _8919_/A _8875_/D vssd1 vssd1 vccd1 vccd1 _8876_/A sky130_fd_sc_hd__or4_4
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7826_ _7761_/X _7821_/Y _7667_/B vssd1 vssd1 vccd1 vccd1 _7826_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_196_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7757_ _9928_/Q vssd1 vssd1 vccd1 vccd1 _8174_/A sky130_fd_sc_hd__inv_2
X_4969_ _4969_/A _4969_/B vssd1 vssd1 vccd1 vccd1 _4969_/Y sky130_fd_sc_hd__nor2_1
XPHY_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7688_ _9926_/Q vssd1 vssd1 vccd1 vccd1 _7901_/A sky130_fd_sc_hd__inv_2
XFILLER_165_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6708_ _6706_/X _6707_/X _6706_/X _6707_/X vssd1 vssd1 vccd1 vccd1 _6716_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9427_ _6571_/Y _6574_/Y _9683_/Q vssd1 vssd1 vccd1 vccd1 _9427_/X sky130_fd_sc_hd__mux2_2
X_6639_ _6760_/A vssd1 vssd1 vccd1 vccd1 _6683_/A sky130_fd_sc_hd__buf_1
XFILLER_192_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9358_ _7062_/A _7618_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9358_/X sky130_fd_sc_hd__mux2_1
X_9289_ _9288_/X _7853_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9289_/X sky130_fd_sc_hd__mux2_1
X_8309_ _7755_/X _9539_/Q _7726_/X _9538_/Q vssd1 vssd1 vccd1 vccd1 _8328_/B sky130_fd_sc_hd__a22o_1
XFILLER_3_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6990_ _6668_/A _6674_/A _6668_/Y vssd1 vssd1 vccd1 vccd1 _6990_/X sky130_fd_sc_hd__a21o_1
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5941_ _9158_/X _5937_/X _9582_/Q _5938_/X vssd1 vssd1 vccd1 vccd1 _9582_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8660_ _8563_/X _8659_/X _8563_/X _8659_/X vssd1 vssd1 vccd1 vccd1 _8660_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_178_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5872_ _9623_/Q vssd1 vssd1 vccd1 vccd1 _5872_/X sky130_fd_sc_hd__buf_2
XFILLER_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8591_ _8591_/A _8591_/B vssd1 vssd1 vccd1 vccd1 _8715_/A sky130_fd_sc_hd__nor2_2
X_4823_ _9908_/Q vssd1 vssd1 vccd1 vccd1 _7665_/A sky130_fd_sc_hd__clkbuf_2
X_7611_ _7602_/A _7602_/B _7603_/B vssd1 vssd1 vccd1 vccd1 _7611_/X sky130_fd_sc_hd__a21bo_1
XFILLER_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4754_ _9525_/Q _9376_/X vssd1 vssd1 vccd1 vccd1 _4754_/X sky130_fd_sc_hd__and2_1
X_7542_ _7540_/X _7541_/X _7540_/X _7541_/X vssd1 vssd1 vccd1 vccd1 _7542_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_193_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7473_ _7473_/A vssd1 vssd1 vccd1 vccd1 _7473_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9212_ _9817_/Q _7642_/Y _9528_/Q vssd1 vssd1 vccd1 vccd1 _9212_/X sky130_fd_sc_hd__mux2_1
X_6424_ _9799_/Q _6537_/B vssd1 vssd1 vccd1 vccd1 _6424_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6355_ _9753_/Q vssd1 vssd1 vccd1 vccd1 _6371_/A sky130_fd_sc_hd__inv_2
XFILLER_115_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9143_ _6145_/X _5035_/A _9148_/S vssd1 vssd1 vccd1 vccd1 _9143_/X sky130_fd_sc_hd__mux2_1
X_6286_ _8036_/A _6142_/A _8038_/A _6141_/A vssd1 vssd1 vccd1 vccd1 _6286_/X sky130_fd_sc_hd__o22a_1
XFILLER_142_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9074_ _6162_/X _5029_/A _9155_/S vssd1 vssd1 vccd1 vccd1 _9074_/X sky130_fd_sc_hd__mux2_1
X_5306_ _9734_/Q _5305_/Y _5240_/A _5305_/A _5224_/X vssd1 vssd1 vccd1 vccd1 _5306_/X
+ sky130_fd_sc_hd__a221o_1
X_8025_ _8025_/A vssd1 vssd1 vccd1 vccd1 _8037_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_102_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5237_ _9732_/Q vssd1 vssd1 vccd1 vccd1 _5238_/B sky130_fd_sc_hd__inv_2
XFILLER_130_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5168_ _5179_/A vssd1 vssd1 vccd1 vccd1 _5168_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5099_ _5115_/A _5099_/B vssd1 vssd1 vccd1 vccd1 _9801_/D sky130_fd_sc_hd__nor2_1
X_8927_ _8927_/A _8927_/B vssd1 vssd1 vccd1 vccd1 _8927_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8858_ _8812_/A _8812_/B _8857_/Y _8812_/Y _8857_/A vssd1 vssd1 vccd1 vccd1 _8859_/B
+ sky130_fd_sc_hd__a32o_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8789_ _8765_/Y _8788_/X _8765_/Y _8788_/X vssd1 vssd1 vccd1 vccd1 _8789_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7809_ _7769_/Y _7805_/Y _7663_/B vssd1 vssd1 vccd1 vccd1 _7809_/Y sky130_fd_sc_hd__o21ai_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6140_ _6140_/A vssd1 vssd1 vccd1 vccd1 _6141_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6071_ _6071_/A vssd1 vssd1 vccd1 vccd1 _6071_/Y sky130_fd_sc_hd__inv_2
X_5022_ _9822_/Q _5019_/X input17/X _5020_/X _5016_/X vssd1 vssd1 vccd1 vccd1 _9822_/D
+ sky130_fd_sc_hd__o221a_1
X_9830_ _9916_/CLK _9830_/D vssd1 vssd1 vccd1 vccd1 _9830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6973_ _6650_/X _6653_/X _6654_/X _6675_/X _6630_/X vssd1 vssd1 vccd1 vccd1 _6973_/X
+ sky130_fd_sc_hd__o221a_1
X_9761_ _9761_/CLK _9761_/D vssd1 vssd1 vccd1 vccd1 _9761_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_19_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8712_ _8773_/C _8766_/B _8712_/C vssd1 vssd1 vccd1 vccd1 _8712_/X sky130_fd_sc_hd__or3_1
X_5924_ _5938_/A vssd1 vssd1 vccd1 vccd1 _5924_/X sky130_fd_sc_hd__buf_2
X_9692_ _9692_/CLK _9692_/D vssd1 vssd1 vccd1 vccd1 _9692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5855_ _9630_/Q vssd1 vssd1 vccd1 vccd1 _8823_/A sky130_fd_sc_hd__buf_2
XFILLER_179_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8643_ _8686_/A _8642_/B _8642_/X vssd1 vssd1 vccd1 vccd1 _8644_/A sky130_fd_sc_hd__a21bo_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4806_ _4830_/A vssd1 vssd1 vccd1 vccd1 _4806_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8574_ _8573_/A _8573_/B _8619_/B vssd1 vssd1 vccd1 vccd1 _8574_/X sky130_fd_sc_hd__a21o_1
XFILLER_194_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5786_ _9659_/Q _5774_/X _5769_/X _7107_/A _5772_/X vssd1 vssd1 vccd1 vccd1 _9659_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_147_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7525_ _7496_/X _7524_/Y _7496_/X _7524_/Y vssd1 vssd1 vccd1 vccd1 _7525_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_21_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7456_ _7355_/X _7370_/X _7355_/X _7370_/X vssd1 vssd1 vccd1 vccd1 _7457_/B sky130_fd_sc_hd__a2bb2o_1
X_6407_ _6407_/A vssd1 vssd1 vccd1 vccd1 _6407_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9126_ _9610_/Q input22/X _9667_/Q vssd1 vssd1 vccd1 vccd1 _9126_/X sky130_fd_sc_hd__mux2_1
X_7387_ _7385_/X _7386_/X _7385_/X _7386_/X vssd1 vssd1 vccd1 vccd1 _7393_/A sky130_fd_sc_hd__a2bb2o_1
X_6338_ _9789_/Q vssd1 vssd1 vccd1 vccd1 _6338_/Y sky130_fd_sc_hd__inv_2
X_6269_ _6268_/A _6268_/B _6268_/X vssd1 vssd1 vccd1 vccd1 _6269_/Y sky130_fd_sc_hd__a21boi_1
X_9057_ _8020_/X _8019_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9057_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8008_ _8008_/A _8008_/B vssd1 vssd1 vccd1 vccd1 _8008_/X sky130_fd_sc_hd__or2_1
XFILLER_84_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5640_ _9680_/Q vssd1 vssd1 vccd1 vccd1 _6596_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5571_ _5482_/X _5539_/X _5482_/X _5539_/X vssd1 vssd1 vccd1 vccd1 _5571_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_191_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8290_ _7728_/X _8212_/Y _8289_/Y vssd1 vssd1 vccd1 vccd1 _8290_/X sky130_fd_sc_hd__o21a_1
XFILLER_144_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7310_ _7311_/A _7385_/B _7313_/C _7379_/A vssd1 vssd1 vccd1 vccd1 _7312_/A sky130_fd_sc_hd__o22a_1
XFILLER_116_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7241_ _7237_/X _7240_/X _7237_/X _7240_/X vssd1 vssd1 vccd1 vccd1 _7241_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_171_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7172_ _7168_/X _7171_/X _7168_/X _7171_/X vssd1 vssd1 vccd1 vccd1 _7172_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_112_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6123_ _9564_/Q _6126_/A _9564_/Q _6126_/A vssd1 vssd1 vccd1 vccd1 _6123_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6054_ _9644_/Q vssd1 vssd1 vccd1 vccd1 _6055_/B sky130_fd_sc_hd__inv_2
XFILLER_58_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5005_ _9833_/Q _5003_/X input29/X _5004_/X _5000_/X vssd1 vssd1 vccd1 vccd1 _9833_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9813_ _9819_/CLK _9813_/D vssd1 vssd1 vccd1 vccd1 _9813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9744_ _9887_/CLK _9744_/D vssd1 vssd1 vccd1 vccd1 _9744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6956_ _6941_/X _6954_/Y _6955_/X vssd1 vssd1 vccd1 vccd1 _6957_/A sky130_fd_sc_hd__a21oi_2
XFILLER_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5907_ _5909_/A _9135_/X vssd1 vssd1 vccd1 vccd1 _9603_/D sky130_fd_sc_hd__and2_1
XFILLER_201_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9675_ _9699_/CLK _9675_/D vssd1 vssd1 vccd1 vccd1 _9675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6887_ _6876_/A _6876_/B _6876_/X vssd1 vssd1 vccd1 vccd1 _6888_/B sky130_fd_sc_hd__a21bo_1
XFILLER_194_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8626_ _8773_/C _8626_/B _8626_/C vssd1 vssd1 vccd1 vccd1 _8626_/X sky130_fd_sc_hd__or3_4
X_5838_ _9638_/Q _5832_/X _5035_/X _5833_/X _5830_/X vssd1 vssd1 vccd1 vccd1 _9638_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_194_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8557_ _8389_/A _8389_/B _8389_/Y vssd1 vssd1 vccd1 vccd1 _8557_/X sky130_fd_sc_hd__a21o_1
X_5769_ _5787_/A vssd1 vssd1 vccd1 vccd1 _5769_/X sky130_fd_sc_hd__buf_1
XFILLER_135_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7508_ _7500_/X _7504_/X _7506_/X _7507_/X vssd1 vssd1 vccd1 vccd1 _7508_/X sky130_fd_sc_hd__o22a_1
XFILLER_175_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8488_ _9689_/Q _8391_/B _8391_/Y vssd1 vssd1 vccd1 vccd1 _8488_/X sky130_fd_sc_hd__a21o_1
XFILLER_190_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7439_ _7294_/X _7372_/Y _7376_/A vssd1 vssd1 vccd1 vccd1 _7439_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_146_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9109_ _6106_/Y _6107_/Y _9896_/Q vssd1 vssd1 vccd1 vccd1 _9109_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6810_ _6795_/X _6796_/X _6808_/X _6809_/X vssd1 vssd1 vccd1 vccd1 _6810_/X sky130_fd_sc_hd__o22a_1
XFILLER_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7790_ _7839_/A vssd1 vssd1 vccd1 vccd1 _7790_/X sky130_fd_sc_hd__buf_4
XFILLER_63_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6741_ _6717_/C _6714_/B _6714_/Y vssd1 vssd1 vccd1 vccd1 _6742_/B sky130_fd_sc_hd__o21ai_1
XFILLER_204_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9460_ _9459_/X _9771_/Q _9481_/S vssd1 vssd1 vccd1 vccd1 _9460_/X sky130_fd_sc_hd__mux2_1
X_6672_ _6672_/A _6672_/B vssd1 vssd1 vccd1 vccd1 _6673_/B sky130_fd_sc_hd__or2_2
XFILLER_176_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5623_ _9701_/Q vssd1 vssd1 vccd1 vccd1 _7637_/A sky130_fd_sc_hd__inv_2
X_8411_ _9698_/Q _6598_/X _8379_/X _8410_/X vssd1 vssd1 vccd1 vccd1 _8411_/X sky130_fd_sc_hd__o22a_2
X_9391_ _9390_/X _9767_/Q _9481_/S vssd1 vssd1 vccd1 vccd1 _9391_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8342_ _9548_/Q vssd1 vssd1 vccd1 vccd1 _8342_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5554_ _5554_/A vssd1 vssd1 vccd1 vccd1 _5554_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8273_ _7666_/A _8234_/Y _8272_/Y vssd1 vssd1 vccd1 vccd1 _8273_/Y sky130_fd_sc_hd__a21oi_1
X_5485_ _5483_/Y _5484_/Y _5483_/Y _5484_/Y vssd1 vssd1 vccd1 vccd1 _5485_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7224_ _7394_/A _7238_/B vssd1 vssd1 vccd1 vccd1 _7224_/X sky130_fd_sc_hd__or2_1
XFILLER_132_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7155_ _7195_/A _9458_/X vssd1 vssd1 vccd1 vccd1 _7155_/X sky130_fd_sc_hd__or2_1
X_6106_ _6103_/X _6105_/X _6103_/X _6105_/X vssd1 vssd1 vccd1 vccd1 _6106_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_86_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7086_ _7086_/A _7086_/B vssd1 vssd1 vccd1 vccd1 _7087_/B sky130_fd_sc_hd__or2_1
X_6037_ _7962_/A _9641_/Q _6026_/A _6028_/Y vssd1 vssd1 vccd1 vccd1 _6037_/X sky130_fd_sc_hd__a22o_1
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7988_ _7988_/A _7993_/B vssd1 vssd1 vccd1 vccd1 _7988_/Y sky130_fd_sc_hd__nor2_1
XPHY_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9727_ _9874_/CLK _9727_/D vssd1 vssd1 vccd1 vccd1 _9727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6939_ _6838_/X _6853_/X _6838_/X _6853_/X vssd1 vssd1 vccd1 vccd1 _6941_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9658_ _9673_/CLK _9658_/D vssd1 vssd1 vccd1 vccd1 _9658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8609_ _8609_/A vssd1 vssd1 vccd1 vccd1 _8702_/C sky130_fd_sc_hd__inv_2
XPHY_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9589_ _9836_/CLK _9589_/D vssd1 vssd1 vccd1 vccd1 _9589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5270_ _5270_/A vssd1 vssd1 vccd1 vccd1 _9743_/D sky130_fd_sc_hd__inv_2
XFILLER_114_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8960_ _8958_/X _8959_/Y _8958_/X _8959_/Y vssd1 vssd1 vccd1 vccd1 _8960_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_209_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7911_ _7911_/A vssd1 vssd1 vccd1 vccd1 _9504_/S sky130_fd_sc_hd__clkinv_8
X_8891_ _8845_/A _8845_/B _8890_/A _8944_/A _8944_/B vssd1 vssd1 vccd1 vccd1 _8891_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_36_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7842_ _7715_/X _7840_/B _7839_/X _7841_/Y vssd1 vssd1 vccd1 vccd1 _7842_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_36_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4985_ _5003_/A vssd1 vssd1 vccd1 vccd1 _4985_/X sky130_fd_sc_hd__clkbuf_2
X_7773_ _7773_/A _7773_/B _7773_/C _7773_/D vssd1 vssd1 vccd1 vccd1 _7773_/X sky130_fd_sc_hd__and4_1
X_6724_ _6720_/X _6723_/X _6720_/X _6723_/X vssd1 vssd1 vccd1 vccd1 _6724_/X sky130_fd_sc_hd__a2bb2o_1
X_9512_ _9844_/Q _9019_/X _7948_/Y _9020_/X _8970_/X _9053_/S vssd1 vssd1 vccd1 vccd1
+ _9512_/X sky130_fd_sc_hd__mux4_2
XPHY_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9443_ _9442_/X _6347_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _9443_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6655_ _6764_/A _9463_/X _6766_/A _6660_/B vssd1 vssd1 vccd1 vccd1 _6656_/A sky130_fd_sc_hd__o22a_1
XFILLER_31_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5606_ _9704_/Q vssd1 vssd1 vccd1 vccd1 _7640_/A sky130_fd_sc_hd__inv_2
X_9374_ _9373_/X _7490_/A _9506_/S vssd1 vssd1 vccd1 vccd1 _9374_/X sky130_fd_sc_hd__mux2_1
X_6586_ _6586_/A vssd1 vssd1 vccd1 vccd1 _6821_/B sky130_fd_sc_hd__buf_1
XFILLER_191_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8325_ _4843_/X _8050_/Y _8320_/Y _8323_/X _8373_/B vssd1 vssd1 vccd1 vccd1 _8325_/Y
+ sky130_fd_sc_hd__o221ai_2
X_5537_ _9385_/X _5487_/X _5581_/A vssd1 vssd1 vccd1 vccd1 _5574_/B sky130_fd_sc_hd__o21ai_1
XFILLER_191_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8256_ _9898_/Q _8254_/X _8255_/X vssd1 vssd1 vccd1 vccd1 _8257_/B sky130_fd_sc_hd__o21ai_1
XFILLER_172_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5468_ _5464_/Y _5467_/X _5464_/Y _5467_/X vssd1 vssd1 vccd1 vccd1 _5549_/A sky130_fd_sc_hd__a2bb2o_1
X_7207_ _7194_/X _7205_/X _7194_/X _7205_/X vssd1 vssd1 vccd1 vccd1 _7207_/X sky130_fd_sc_hd__a2bb2o_1
X_8187_ _8187_/A _8187_/B vssd1 vssd1 vccd1 vccd1 _8187_/Y sky130_fd_sc_hd__nor2_1
X_5399_ _5396_/Y _5397_/Y _5398_/Y vssd1 vssd1 vccd1 vccd1 _5399_/X sky130_fd_sc_hd__o21a_1
XFILLER_98_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7138_ _7522_/A _7490_/B _7494_/A _7169_/B vssd1 vssd1 vccd1 vccd1 _7138_/X sky130_fd_sc_hd__o22a_1
XFILLER_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7069_ _7069_/A _7069_/B vssd1 vssd1 vccd1 vccd1 _7070_/B sky130_fd_sc_hd__nand2_1
XFILLER_100_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 io_wb_dat_i[12] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_4
XFILLER_182_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4770_ _7684_/A vssd1 vssd1 vccd1 vccd1 _4770_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6440_ _9792_/Q _6528_/B vssd1 vssd1 vccd1 vccd1 _6463_/A sky130_fd_sc_hd__nor2_1
XFILLER_173_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6371_ _6371_/A _6371_/B vssd1 vssd1 vccd1 vccd1 _6372_/B sky130_fd_sc_hd__nand2_1
XFILLER_173_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8110_ _9544_/Q _8072_/B _8073_/B vssd1 vssd1 vccd1 vccd1 _8110_/X sky130_fd_sc_hd__a21bo_1
X_5322_ _9722_/Q vssd1 vssd1 vccd1 vccd1 _5329_/A sky130_fd_sc_hd__inv_2
X_9090_ _9089_/X _7858_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9090_/X sky130_fd_sc_hd__mux2_1
X_8041_ _9441_/X _8045_/B vssd1 vssd1 vccd1 vccd1 _8041_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5253_ _5271_/A vssd1 vssd1 vccd1 vccd1 _5253_/Y sky130_fd_sc_hd__inv_2
X_5184_ _6351_/A _5178_/X input25/X _5179_/X _5175_/X vssd1 vssd1 vccd1 vccd1 _9766_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_87_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8943_ _8922_/X _8923_/X _8881_/X _8924_/X vssd1 vssd1 vccd1 vccd1 _8943_/X sky130_fd_sc_hd__o22a_1
X_8874_ _8863_/X _8873_/X _8863_/X _8873_/X vssd1 vssd1 vccd1 vccd1 _8874_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7825_ _7696_/X _7823_/B _7781_/A _7824_/Y vssd1 vssd1 vccd1 vccd1 _7825_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_24_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7756_ _9927_/Q vssd1 vssd1 vccd1 vccd1 _7906_/A sky130_fd_sc_hd__inv_2
XFILLER_149_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4968_ _5026_/A vssd1 vssd1 vccd1 vccd1 _4968_/Y sky130_fd_sc_hd__inv_2
XPHY_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7687_ _8257_/A vssd1 vssd1 vccd1 vccd1 _8134_/A sky130_fd_sc_hd__clkbuf_2
X_6707_ _6707_/A _6721_/B vssd1 vssd1 vccd1 vccd1 _6707_/X sky130_fd_sc_hd__or2_1
X_4899_ _5586_/A vssd1 vssd1 vccd1 vccd1 _5787_/A sky130_fd_sc_hd__buf_2
XPHY_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6638_ _6634_/X _6637_/X _6634_/X _6637_/X vssd1 vssd1 vccd1 vccd1 _6646_/A sky130_fd_sc_hd__a2bb2o_1
X_9426_ _6569_/Y _6570_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9426_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9357_ _7623_/X _7586_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9357_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6569_ _6569_/A vssd1 vssd1 vccd1 vccd1 _6569_/Y sky130_fd_sc_hd__inv_2
X_8308_ _9540_/Q vssd1 vssd1 vccd1 vccd1 _8308_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9288_ _9766_/Q _9287_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9288_/X sky130_fd_sc_hd__mux2_1
X_8239_ _9757_/Q _8243_/A vssd1 vssd1 vccd1 vccd1 _8240_/B sky130_fd_sc_hd__or2_2
XFILLER_105_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5940_ _9159_/X _5937_/X _9583_/Q _5938_/X vssd1 vssd1 vccd1 vccd1 _9583_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7610_ _7079_/A _7079_/B _7080_/B vssd1 vssd1 vccd1 vccd1 _7610_/X sky130_fd_sc_hd__a21bo_1
X_5871_ _7210_/A _5865_/X _5032_/X _5866_/X _5867_/X vssd1 vssd1 vccd1 vccd1 _9624_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8590_ _8589_/A _8589_/B _8633_/A vssd1 vssd1 vccd1 vccd1 _8591_/B sky130_fd_sc_hd__a21o_1
X_4822_ _4834_/A vssd1 vssd1 vccd1 vccd1 _4822_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4753_ _4753_/A vssd1 vssd1 vccd1 vccd1 _4753_/Y sky130_fd_sc_hd__inv_2
X_7541_ _7190_/A _7190_/B _7191_/B vssd1 vssd1 vccd1 vccd1 _7541_/X sky130_fd_sc_hd__a21bo_1
XFILLER_159_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7472_ _7457_/X _7470_/Y _7471_/X vssd1 vssd1 vccd1 vccd1 _7473_/A sky130_fd_sc_hd__a21oi_2
X_9211_ _9816_/Q _7640_/Y _9528_/Q vssd1 vssd1 vccd1 vccd1 _9211_/X sky130_fd_sc_hd__mux2_1
X_6423_ _6423_/A vssd1 vssd1 vccd1 vccd1 _6537_/B sky130_fd_sc_hd__inv_2
XFILLER_174_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6354_ _9779_/Q vssd1 vssd1 vccd1 vccd1 _6354_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9142_ _6124_/X _5039_/A _9155_/S vssd1 vssd1 vccd1 vccd1 _9142_/X sky130_fd_sc_hd__mux2_1
X_6285_ _6285_/A _6275_/X vssd1 vssd1 vccd1 vccd1 _6285_/X sky130_fd_sc_hd__or2b_1
X_9073_ _6121_/Y _5041_/A _9155_/S vssd1 vssd1 vccd1 vccd1 _9073_/X sky130_fd_sc_hd__mux2_1
X_5305_ _5305_/A vssd1 vssd1 vccd1 vccd1 _5305_/Y sky130_fd_sc_hd__inv_2
X_8024_ _8024_/A _8033_/B vssd1 vssd1 vccd1 vccd1 _8024_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5236_ _9733_/Q vssd1 vssd1 vccd1 vccd1 _5238_/A sky130_fd_sc_hd__inv_2
XFILLER_130_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5167_ _5178_/A vssd1 vssd1 vccd1 vccd1 _5167_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5098_ _5084_/X _6318_/C _5096_/Y _5097_/X vssd1 vssd1 vccd1 vccd1 _5099_/B sky130_fd_sc_hd__o22a_1
XFILLER_83_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8926_ _8899_/X _8925_/X _8899_/X _8925_/X vssd1 vssd1 vccd1 vccd1 _8926_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8857_ _8857_/A vssd1 vssd1 vccd1 vccd1 _8857_/Y sky130_fd_sc_hd__inv_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8788_ _8786_/X _8788_/B vssd1 vssd1 vccd1 vccd1 _8788_/X sky130_fd_sc_hd__and2b_1
X_7808_ _7807_/A _7807_/B _7810_/B _7839_/A vssd1 vssd1 vccd1 vccd1 _7808_/Y sky130_fd_sc_hd__a211oi_4
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7739_ _9926_/Q _6343_/Y _7738_/X _6351_/A vssd1 vssd1 vccd1 vccd1 _7739_/X sky130_fd_sc_hd__o22a_1
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9409_ _9408_/X _6331_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _9409_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6070_ _7981_/A _9644_/Q _6056_/B _6061_/X vssd1 vssd1 vccd1 vccd1 _6071_/A sky130_fd_sc_hd__o22a_1
X_5021_ _9823_/Q _5019_/X input18/X _5020_/X _5016_/X vssd1 vssd1 vccd1 vccd1 _9823_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9760_ _9909_/CLK _9760_/D vssd1 vssd1 vccd1 vccd1 _9760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8711_ _8668_/Y _8671_/X _8672_/X _8673_/X vssd1 vssd1 vccd1 vccd1 _8711_/X sky130_fd_sc_hd__o22a_1
X_6972_ _9617_/Q _6691_/B _6970_/A _6970_/Y _6971_/X vssd1 vssd1 vccd1 vccd1 _6972_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_65_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9691_ _9692_/CLK _9691_/D vssd1 vssd1 vccd1 vccd1 _9691_/Q sky130_fd_sc_hd__dfxtp_1
X_5923_ _5959_/A vssd1 vssd1 vccd1 vccd1 _5938_/A sky130_fd_sc_hd__buf_4
XFILLER_34_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5854_ _5852_/X _5847_/X _4978_/X _5848_/X _5853_/X vssd1 vssd1 vccd1 vccd1 _9631_/D
+ sky130_fd_sc_hd__o221a_1
X_8642_ _8686_/A _8642_/B vssd1 vssd1 vccd1 vccd1 _8642_/X sky130_fd_sc_hd__or2_1
XFILLER_110_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8573_ _8573_/A _8573_/B vssd1 vssd1 vccd1 vccd1 _8619_/B sky130_fd_sc_hd__nor2_2
XFILLER_194_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4805_ _9091_/X _4796_/X _7673_/A _4799_/X _4791_/X vssd1 vssd1 vccd1 vccd1 _9916_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5785_ _5785_/A vssd1 vssd1 vccd1 vccd1 _7107_/A sky130_fd_sc_hd__inv_2
X_7524_ _7520_/X _7523_/X _7520_/X _7523_/X vssd1 vssd1 vccd1 vccd1 _7524_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_21_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7455_ _7420_/A _7420_/B _7442_/B vssd1 vssd1 vccd1 vccd1 _7457_/A sky130_fd_sc_hd__a21o_1
X_6406_ _5162_/X _6393_/B _8199_/A vssd1 vssd1 vccd1 vccd1 _6546_/B sky130_fd_sc_hd__a21boi_2
X_7386_ _7386_/A _7398_/B vssd1 vssd1 vccd1 vccd1 _7386_/X sky130_fd_sc_hd__or2_1
XFILLER_150_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6337_ _6337_/A vssd1 vssd1 vccd1 vccd1 _6337_/Y sky130_fd_sc_hd__inv_2
X_9125_ _9609_/Q input21/X _9667_/Q vssd1 vssd1 vccd1 vccd1 _9125_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6268_ _6268_/A _6268_/B vssd1 vssd1 vccd1 vccd1 _6268_/X sky130_fd_sc_hd__or2_2
X_9056_ _8018_/Y _8017_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9056_/X sky130_fd_sc_hd__mux2_1
X_5219_ _5039_/X _5151_/X _5218_/X _5152_/X _5214_/X vssd1 vssd1 vccd1 vccd1 _9749_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8007_ _9409_/X _8022_/B vssd1 vssd1 vccd1 vccd1 _8007_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6199_ _6199_/A vssd1 vssd1 vccd1 vccd1 _6221_/A sky130_fd_sc_hd__inv_2
XFILLER_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8909_ _9419_/X vssd1 vssd1 vccd1 vccd1 _8909_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9889_ _9893_/CLK _9889_/D vssd1 vssd1 vccd1 vccd1 _9889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5570_ _5787_/A vssd1 vssd1 vccd1 vccd1 _5570_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7240_ _7490_/A _7283_/B _7240_/C vssd1 vssd1 vccd1 vccd1 _7240_/X sky130_fd_sc_hd__or3_1
XFILLER_7_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7171_ _7491_/A _7494_/B _7171_/C vssd1 vssd1 vccd1 vccd1 _7171_/X sky130_fd_sc_hd__or3_1
XFILLER_124_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6122_ _5969_/Y _9521_/Q _9518_/D _5972_/Y vssd1 vssd1 vccd1 vccd1 _6126_/A sky130_fd_sc_hd__o22a_2
XFILLER_112_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6053_ _7981_/A _9644_/Q vssd1 vssd1 vccd1 vccd1 _6056_/A sky130_fd_sc_hd__nor2_1
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5004_ _5004_/A vssd1 vssd1 vccd1 vccd1 _5004_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9812_ _9819_/CLK _9812_/D vssd1 vssd1 vccd1 vccd1 _9812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9743_ _9893_/CLK _9743_/D vssd1 vssd1 vccd1 vccd1 _9743_/Q sky130_fd_sc_hd__dfxtp_1
X_6955_ _6713_/C _6936_/X _6713_/C _6936_/X vssd1 vssd1 vccd1 vccd1 _6955_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9674_ _9699_/CLK _9674_/D vssd1 vssd1 vccd1 vccd1 _9674_/Q sky130_fd_sc_hd__dfxtp_1
X_5906_ _5909_/A _9136_/X vssd1 vssd1 vccd1 vccd1 _9604_/D sky130_fd_sc_hd__and2_1
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8625_ _8773_/A _8625_/B vssd1 vssd1 vccd1 vccd1 _8766_/C sky130_fd_sc_hd__or2_2
X_6886_ _6886_/A _6867_/X vssd1 vssd1 vccd1 vccd1 _6888_/A sky130_fd_sc_hd__or2b_1
XFILLER_194_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5837_ _4978_/X _5818_/X _9639_/Q _5819_/X _5214_/X vssd1 vssd1 vccd1 vccd1 _9639_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8556_ _8555_/A _8555_/B _8599_/A vssd1 vssd1 vccd1 vccd1 _8556_/X sky130_fd_sc_hd__a21bo_1
X_5768_ _9664_/Q _5697_/X _5570_/X _7121_/A _5698_/X vssd1 vssd1 vccd1 vccd1 _9664_/D
+ sky130_fd_sc_hd__o221a_1
X_8487_ _8486_/A _8486_/B _8522_/A vssd1 vssd1 vccd1 vccd1 _8487_/X sky130_fd_sc_hd__a21bo_1
X_7507_ _7500_/X _7504_/X _7500_/X _7504_/X vssd1 vssd1 vccd1 vccd1 _7507_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_147_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5699_ _6571_/A _5697_/X _9096_/X _5692_/X _5698_/X vssd1 vssd1 vccd1 vccd1 _9669_/D
+ sky130_fd_sc_hd__o221a_1
X_7438_ _7434_/X _7435_/X _7434_/X _7435_/X vssd1 vssd1 vccd1 vccd1 _7438_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_190_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7369_ _7361_/X _7364_/X _7367_/X _7368_/X vssd1 vssd1 vccd1 vccd1 _7369_/X sky130_fd_sc_hd__o22a_1
X_9108_ _6097_/X _6099_/X _9896_/Q vssd1 vssd1 vccd1 vccd1 _9108_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9039_ _7993_/Y _9606_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9039_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6740_ _6728_/A _6728_/B _6910_/A vssd1 vssd1 vccd1 vccd1 _6743_/A sky130_fd_sc_hd__a21o_1
XFILLER_63_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6671_ _6647_/C _6644_/B _6644_/Y vssd1 vssd1 vccd1 vccd1 _6672_/B sky130_fd_sc_hd__o21ai_1
XFILLER_31_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5622_ _5626_/A _5622_/B vssd1 vssd1 vccd1 vccd1 _5622_/X sky130_fd_sc_hd__and2_1
X_8410_ _9697_/Q _6591_/Y _8381_/Y _8409_/X vssd1 vssd1 vccd1 vccd1 _8410_/X sky130_fd_sc_hd__o22a_1
X_9390_ _9799_/Q _9916_/Q _9480_/S vssd1 vssd1 vccd1 vccd1 _9390_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8341_ _7743_/X _9545_/Q _7728_/X _9552_/Q vssd1 vssd1 vccd1 vccd1 _8346_/B sky130_fd_sc_hd__a22o_1
X_5553_ _5692_/A vssd1 vssd1 vccd1 vccd1 _5553_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8272_ _7823_/A _8241_/X _8271_/X vssd1 vssd1 vccd1 vccd1 _8272_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5484_ _5418_/A _5418_/B _5418_/Y vssd1 vssd1 vccd1 vccd1 _5484_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_172_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7223_ _7223_/A _9469_/X vssd1 vssd1 vccd1 vccd1 _7223_/X sky130_fd_sc_hd__or2_1
XFILLER_98_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7154_ _7160_/A vssd1 vssd1 vccd1 vccd1 _7195_/A sky130_fd_sc_hd__buf_1
XFILLER_112_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6105_ _6088_/X _6095_/A _6104_/X vssd1 vssd1 vccd1 vccd1 _6105_/X sky130_fd_sc_hd__o21ba_1
XFILLER_140_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7085_ _7085_/A _7085_/B vssd1 vssd1 vccd1 vccd1 _7086_/B sky130_fd_sc_hd__or2_1
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6036_ _6036_/A vssd1 vssd1 vccd1 vccd1 _6036_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7987_ _9375_/X _7987_/B vssd1 vssd1 vccd1 vccd1 _7987_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9726_ _9874_/CLK _9726_/D vssd1 vssd1 vccd1 vccd1 _9726_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6938_ _6933_/X _6937_/X _6933_/X _6937_/X vssd1 vssd1 vccd1 vccd1 _6938_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9657_ _9673_/CLK _9657_/D vssd1 vssd1 vccd1 vccd1 _9657_/Q sky130_fd_sc_hd__dfxtp_1
X_6869_ _6877_/A _6881_/B vssd1 vssd1 vccd1 vccd1 _6869_/X sky130_fd_sc_hd__or2_1
XFILLER_22_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8608_ _8821_/A _9457_/X vssd1 vssd1 vccd1 vccd1 _8609_/A sky130_fd_sc_hd__or2_2
X_9588_ _9836_/CLK _9588_/D vssd1 vssd1 vccd1 vccd1 _9588_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8539_ _8610_/C _8538_/B _8573_/A vssd1 vssd1 vccd1 vccd1 _8539_/X sky130_fd_sc_hd__a21bo_1
XFILLER_157_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7910_ _8301_/A _7909_/Y _8174_/A _7909_/A _7785_/X vssd1 vssd1 vccd1 vccd1 _7910_/X
+ sky130_fd_sc_hd__o221a_1
X_8890_ _8890_/A vssd1 vssd1 vccd1 vccd1 _8944_/B sky130_fd_sc_hd__inv_2
X_7841_ _7844_/B vssd1 vssd1 vccd1 vccd1 _7841_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7772_ _7772_/A _7772_/B _7772_/C _7772_/D vssd1 vssd1 vccd1 vccd1 _7773_/D sky130_fd_sc_hd__and4_1
X_4984_ _5028_/A vssd1 vssd1 vccd1 vccd1 _5003_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6723_ _7005_/A _6766_/B _6723_/C vssd1 vssd1 vccd1 vccd1 _6723_/X sky130_fd_sc_hd__or3_1
X_9511_ _9528_/Q _9016_/X _7942_/Y _9017_/X _8970_/X _9053_/S vssd1 vssd1 vccd1 vccd1
+ _9511_/X sky130_fd_sc_hd__mux4_2
XFILLER_189_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9442_ _6317_/D _7709_/X _9480_/S vssd1 vssd1 vccd1 vccd1 _9442_/X sky130_fd_sc_hd__mux2_1
X_6654_ _6650_/X _6653_/X _6650_/X _6653_/X vssd1 vssd1 vccd1 vccd1 _6654_/X sky130_fd_sc_hd__a2bb2o_1
X_5605_ _5605_/A _5605_/B vssd1 vssd1 vccd1 vccd1 _5605_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9373_ _9372_/X _8955_/A _9505_/S vssd1 vssd1 vccd1 vccd1 _9373_/X sky130_fd_sc_hd__mux2_1
X_6585_ _9613_/Q vssd1 vssd1 vccd1 vccd1 _6586_/A sky130_fd_sc_hd__inv_2
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8324_ _8324_/A _8324_/B vssd1 vssd1 vccd1 vccd1 _8373_/B sky130_fd_sc_hd__or2_1
X_5536_ _5582_/A _5582_/B vssd1 vssd1 vccd1 vccd1 _5581_/A sky130_fd_sc_hd__nand2_1
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8255_ _8187_/A _8187_/B _9898_/Q _8254_/X _8187_/Y vssd1 vssd1 vccd1 vccd1 _8255_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5467_ _5467_/A _5467_/B vssd1 vssd1 vccd1 vccd1 _5467_/X sky130_fd_sc_hd__and2_1
X_7206_ _7147_/A _7147_/B _7147_/Y vssd1 vssd1 vccd1 vccd1 _7206_/X sky130_fd_sc_hd__a21o_1
X_8186_ _8186_/A _9748_/Q vssd1 vssd1 vccd1 vccd1 _8187_/B sky130_fd_sc_hd__nor2_2
X_5398_ _9718_/Q vssd1 vssd1 vccd1 vccd1 _5398_/Y sky130_fd_sc_hd__inv_2
X_7137_ _7169_/B vssd1 vssd1 vccd1 vccd1 _7137_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7068_ _7068_/A vssd1 vssd1 vccd1 vccd1 _7069_/B sky130_fd_sc_hd__inv_2
XFILLER_100_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6019_ _6019_/A vssd1 vssd1 vccd1 vccd1 _6019_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9709_ _9828_/CLK _9709_/D vssd1 vssd1 vccd1 vccd1 _9709_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6370_ _4960_/X _8191_/A _6359_/Y _6369_/X vssd1 vssd1 vccd1 vccd1 _6371_/B sky130_fd_sc_hd__o22a_1
XFILLER_127_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5321_ _9723_/Q vssd1 vssd1 vccd1 vccd1 _5330_/A sky130_fd_sc_hd__inv_2
X_8040_ _8040_/A _8044_/B vssd1 vssd1 vccd1 vccd1 _8040_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5252_ _9747_/Q vssd1 vssd1 vccd1 vccd1 _5252_/Y sky130_fd_sc_hd__inv_2
X_5183_ _9766_/Q vssd1 vssd1 vccd1 vccd1 _6351_/A sky130_fd_sc_hd__buf_2
XFILLER_68_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8942_ _8942_/A _8942_/B vssd1 vssd1 vccd1 vccd1 _8942_/Y sky130_fd_sc_hd__nor2_1
X_8873_ _8903_/A _8833_/B _8872_/Y _8833_/Y _8872_/A vssd1 vssd1 vccd1 vccd1 _8873_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_64_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7824_ _7827_/B vssd1 vssd1 vccd1 vccd1 _7824_/Y sky130_fd_sc_hd__inv_2
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4967_ _5032_/A vssd1 vssd1 vccd1 vccd1 _4969_/B sky130_fd_sc_hd__inv_2
X_7755_ _7819_/A vssd1 vssd1 vccd1 vccd1 _7755_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7686_ _9899_/Q vssd1 vssd1 vccd1 vccd1 _8257_/A sky130_fd_sc_hd__inv_2
XFILLER_149_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4898_ _5339_/A vssd1 vssd1 vccd1 vccd1 _5586_/A sky130_fd_sc_hd__clkbuf_4
X_6706_ _6706_/A _6760_/B vssd1 vssd1 vccd1 vccd1 _6706_/X sky130_fd_sc_hd__or2_1
XFILLER_177_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6637_ _6760_/A _9462_/X vssd1 vssd1 vccd1 vccd1 _6637_/X sky130_fd_sc_hd__or2_1
X_9425_ _6567_/Y _6568_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9425_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6568_ _8394_/B _6554_/B _6565_/Y vssd1 vssd1 vccd1 vccd1 _6568_/X sky130_fd_sc_hd__a21o_1
X_9356_ _7059_/A _7612_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9356_/X sky130_fd_sc_hd__mux2_1
X_5519_ _9490_/X _5510_/X _9490_/X _5510_/X vssd1 vssd1 vccd1 vccd1 _5622_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_145_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8307_ _4816_/X _8305_/Y _7666_/A _8306_/Y vssd1 vssd1 vccd1 vccd1 _8328_/C sky130_fd_sc_hd__a22o_1
XFILLER_3_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6499_ _6499_/A vssd1 vssd1 vccd1 vccd1 _6499_/Y sky130_fd_sc_hd__inv_2
X_9287_ _7851_/Y _9766_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9287_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8238_ _9756_/Q _8238_/B vssd1 vssd1 vccd1 vccd1 _8243_/A sky130_fd_sc_hd__or2_1
XFILLER_105_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8169_ _4775_/X _8095_/Y _4780_/X _8096_/Y _8168_/X vssd1 vssd1 vccd1 vccd1 _8169_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_47_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5870_ _9624_/Q vssd1 vssd1 vccd1 vccd1 _7210_/A sky130_fd_sc_hd__buf_2
X_4821_ _9274_/X _4809_/X _4820_/X _4810_/X _4817_/X vssd1 vssd1 vccd1 vccd1 _9909_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4752_ _9282_/S _9525_/D vssd1 vssd1 vccd1 vccd1 _4753_/A sky130_fd_sc_hd__or2b_2
X_7540_ _7474_/X _7475_/X _7474_/X _7475_/X vssd1 vssd1 vccd1 vccd1 _7540_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_147_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7471_ _7230_/C _7452_/X _7230_/C _7452_/X vssd1 vssd1 vccd1 vccd1 _7471_/X sky130_fd_sc_hd__a2bb2o_1
X_9210_ _9815_/Q _7639_/Y _9528_/Q vssd1 vssd1 vccd1 vccd1 _9210_/X sky130_fd_sc_hd__mux2_1
X_6422_ _5181_/X _8219_/A _8215_/A vssd1 vssd1 vccd1 vccd1 _6423_/A sky130_fd_sc_hd__a21bo_1
XFILLER_146_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9141_ _9879_/Q _9895_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9141_/X sky130_fd_sc_hd__mux2_1
X_6353_ _6353_/A vssd1 vssd1 vccd1 vccd1 _6353_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6284_ _9591_/Q _6171_/A _8040_/A _6142_/A vssd1 vssd1 vccd1 vccd1 _6288_/A sky130_fd_sc_hd__a22o_1
XFILLER_142_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9072_ _9876_/Q _9892_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9072_/X sky130_fd_sc_hd__mux2_1
X_5304_ _5304_/A vssd1 vssd1 vccd1 vccd1 _9735_/D sky130_fd_sc_hd__inv_2
X_8023_ _8046_/B vssd1 vssd1 vccd1 vccd1 _8033_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_142_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5235_ _9734_/Q vssd1 vssd1 vccd1 vccd1 _5240_/A sky130_fd_sc_hd__inv_2
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5166_ _8205_/A _5155_/X input34/X _5157_/X _5165_/X vssd1 vssd1 vccd1 vccd1 _9774_/D
+ sky130_fd_sc_hd__o221a_1
X_5097_ _5097_/A vssd1 vssd1 vccd1 vccd1 _5097_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_204_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8925_ _8881_/X _8924_/X _8881_/X _8924_/X vssd1 vssd1 vccd1 vccd1 _8925_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8856_ _8854_/Y _8895_/B _8854_/Y _8895_/B vssd1 vssd1 vccd1 vccd1 _8857_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8787_ _8787_/A _8787_/B vssd1 vssd1 vccd1 vccd1 _8788_/B sky130_fd_sc_hd__or2_1
X_7807_ _7807_/A _7807_/B vssd1 vssd1 vccd1 vccd1 _7810_/B sky130_fd_sc_hd__nor2_4
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5999_ _9850_/Q _5985_/Y _5989_/X vssd1 vssd1 vccd1 vccd1 _5999_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_197_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7738_ _7738_/A vssd1 vssd1 vccd1 vccd1 _7738_/X sky130_fd_sc_hd__buf_2
XFILLER_184_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9408_ _6330_/Y _7713_/X _9480_/S vssd1 vssd1 vccd1 vccd1 _9408_/X sky130_fd_sc_hd__mux2_1
X_7669_ _9912_/Q _7669_/B vssd1 vssd1 vccd1 vccd1 _7837_/A sky130_fd_sc_hd__or2_1
XFILLER_20_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9339_ _7056_/A _7606_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9339_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5020_ _5030_/A vssd1 vssd1 vccd1 vccd1 _5020_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8710_ _8708_/X _8709_/X _8708_/X _8709_/X vssd1 vssd1 vccd1 vccd1 _8710_/X sky130_fd_sc_hd__a2bb2o_1
X_6971_ _6971_/A _6971_/B vssd1 vssd1 vccd1 vccd1 _6971_/X sky130_fd_sc_hd__or2_1
XFILLER_206_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9690_ _9692_/CLK _9690_/D vssd1 vssd1 vccd1 vccd1 _9690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5922_ _5958_/A vssd1 vssd1 vccd1 vccd1 _5959_/A sky130_fd_sc_hd__inv_2
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8641_ _8593_/Y _8596_/Y _8639_/X _8640_/Y vssd1 vssd1 vccd1 vccd1 _8642_/B sky130_fd_sc_hd__o31ai_4
X_5853_ _5891_/A vssd1 vssd1 vccd1 vccd1 _5853_/X sky130_fd_sc_hd__buf_1
XFILLER_80_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8572_ _8571_/A _8571_/B _8619_/A vssd1 vssd1 vccd1 vccd1 _8573_/B sky130_fd_sc_hd__a21o_1
XFILLER_179_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4804_ _9916_/Q vssd1 vssd1 vccd1 vccd1 _7673_/A sky130_fd_sc_hd__buf_1
X_5784_ _5730_/X _5750_/X _5730_/X _5750_/X vssd1 vssd1 vccd1 vccd1 _5785_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_166_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7523_ _7521_/X _7522_/X _7521_/X _7522_/X vssd1 vssd1 vccd1 vccd1 _7523_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7454_ _7449_/X _7453_/X _7449_/X _7453_/X vssd1 vssd1 vccd1 vccd1 _7454_/X sky130_fd_sc_hd__a2bb2o_1
X_6405_ _6405_/A vssd1 vssd1 vccd1 vccd1 _6548_/B sky130_fd_sc_hd__inv_2
XFILLER_174_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7385_ _7385_/A _7385_/B vssd1 vssd1 vccd1 vccd1 _7385_/X sky130_fd_sc_hd__or2_1
XFILLER_162_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6336_ _9790_/Q vssd1 vssd1 vccd1 vccd1 _6453_/A sky130_fd_sc_hd__inv_2
X_9124_ _9608_/Q input20/X _9667_/Q vssd1 vssd1 vccd1 vccd1 _9124_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9055_ _8016_/Y _8015_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9055_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6267_ _6247_/A _6265_/X _6247_/B _6266_/X vssd1 vssd1 vccd1 vccd1 _6268_/B sky130_fd_sc_hd__o211a_1
XFILLER_130_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5218_ _9749_/Q vssd1 vssd1 vccd1 vccd1 _5218_/X sky130_fd_sc_hd__buf_2
X_8006_ _8045_/B vssd1 vssd1 vccd1 vccd1 _8022_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_103_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6198_ _7997_/A _6201_/A _9575_/Q _6166_/A vssd1 vssd1 vccd1 vccd1 _6199_/A sky130_fd_sc_hd__o22a_1
XFILLER_57_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5149_ _5179_/A vssd1 vssd1 vccd1 vccd1 _5178_/A sky130_fd_sc_hd__inv_2
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8908_ _8942_/B vssd1 vssd1 vccd1 vccd1 _8908_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9888_ _9888_/CLK _9888_/D vssd1 vssd1 vccd1 vccd1 _9888_/Q sky130_fd_sc_hd__dfxtp_1
X_8839_ _8837_/X _8838_/X _8837_/X _8838_/X vssd1 vssd1 vccd1 vccd1 _8840_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7170_ _7170_/A vssd1 vssd1 vccd1 vccd1 _7171_/C sky130_fd_sc_hd__inv_2
X_6121_ _9563_/Q vssd1 vssd1 vccd1 vccd1 _6121_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6052_ _9857_/Q vssd1 vssd1 vccd1 vccd1 _7981_/A sky130_fd_sc_hd__inv_2
XFILLER_39_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5003_ _5003_/A vssd1 vssd1 vccd1 vccd1 _5003_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9811_ _9928_/CLK _9811_/D vssd1 vssd1 vccd1 vccd1 _9811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9742_ _9893_/CLK _9742_/D vssd1 vssd1 vccd1 vccd1 _9742_/Q sky130_fd_sc_hd__dfxtp_1
X_6954_ _6954_/A _6954_/B vssd1 vssd1 vccd1 vccd1 _6954_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9673_ _9673_/CLK _9673_/D vssd1 vssd1 vccd1 vccd1 _9673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5905_ _5909_/A _9137_/X vssd1 vssd1 vccd1 vccd1 _9605_/D sky130_fd_sc_hd__and2_1
X_8624_ _8623_/A _8623_/B _8709_/A vssd1 vssd1 vccd1 vccd1 _8624_/X sky130_fd_sc_hd__a21bo_1
X_6885_ _6867_/A _6867_/B _6867_/C _6867_/D vssd1 vssd1 vccd1 vccd1 _6886_/A sky130_fd_sc_hd__o22a_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5836_ _9640_/Q _5832_/X _5032_/X _5833_/X _5830_/X vssd1 vssd1 vccd1 vccd1 _9640_/D
+ sky130_fd_sc_hd__o221a_1
X_8555_ _8555_/A _8555_/B vssd1 vssd1 vccd1 vccd1 _8599_/A sky130_fd_sc_hd__or2_1
X_5767_ _5755_/X _5766_/X _5755_/X _5766_/X vssd1 vssd1 vccd1 vccd1 _7121_/A sky130_fd_sc_hd__o2bb2a_2
XFILLER_194_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8486_ _8486_/A _8486_/B vssd1 vssd1 vccd1 vccd1 _8522_/A sky130_fd_sc_hd__or2_2
XFILLER_135_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5698_ _5772_/A vssd1 vssd1 vccd1 vccd1 _5698_/X sky130_fd_sc_hd__buf_2
X_7506_ _7506_/A _7506_/B vssd1 vssd1 vccd1 vccd1 _7506_/X sky130_fd_sc_hd__or2_1
XFILLER_135_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7437_ _7477_/A _7477_/B vssd1 vssd1 vccd1 vccd1 _7437_/X sky130_fd_sc_hd__and2_1
XFILLER_146_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7368_ _7361_/X _7364_/X _7361_/X _7364_/X vssd1 vssd1 vccd1 vccd1 _7368_/X sky130_fd_sc_hd__a2bb2o_1
X_6319_ _4960_/X _6309_/Y _6316_/X _6317_/X _6318_/X vssd1 vssd1 vccd1 vccd1 _6319_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9107_ _6089_/Y _6090_/Y _9896_/Q vssd1 vssd1 vccd1 vccd1 _9107_/X sky130_fd_sc_hd__mux2_1
X_7299_ _7299_/A vssd1 vssd1 vccd1 vccd1 _7372_/A sky130_fd_sc_hd__inv_2
XFILLER_130_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9038_ _7989_/Y _9037_/X _9038_/S vssd1 vssd1 vccd1 vccd1 _9038_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_1_clock clkbuf_1_1_1_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6670_ _6658_/A _6658_/B _6991_/A vssd1 vssd1 vccd1 vccd1 _6673_/A sky130_fd_sc_hd__a21o_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5621_ _5621_/A vssd1 vssd1 vccd1 vccd1 _5621_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8340_ _8340_/A _8340_/B _8340_/C _8339_/X vssd1 vssd1 vccd1 vccd1 _8346_/A sky130_fd_sc_hd__or4b_4
X_5552_ _9715_/Q _4897_/X _5910_/A _5551_/X vssd1 vssd1 vccd1 vccd1 _9715_/D sky130_fd_sc_hd__o211a_1
XFILLER_191_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8271_ _7823_/A _8241_/X _7819_/A _8242_/X _8270_/X vssd1 vssd1 vccd1 vccd1 _8271_/X
+ sky130_fd_sc_hd__o221a_1
X_5483_ _5483_/A vssd1 vssd1 vccd1 vccd1 _5483_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7222_ _7247_/A _7222_/B _7400_/A _7247_/B vssd1 vssd1 vccd1 vccd1 _7222_/X sky130_fd_sc_hd__or4_4
XFILLER_144_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7153_ _7178_/A _7522_/B _7265_/A _7178_/B vssd1 vssd1 vccd1 vccd1 _7153_/X sky130_fd_sc_hd__or4_4
X_6104_ _7999_/A _9648_/Q _6095_/B _6098_/X vssd1 vssd1 vccd1 vccd1 _6104_/X sky130_fd_sc_hd__o22a_1
XFILLER_86_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7084_ _7084_/A _7084_/B vssd1 vssd1 vccd1 vccd1 _7085_/B sky130_fd_sc_hd__or2_1
X_6035_ _9855_/Q _6034_/B _6034_/Y vssd1 vssd1 vccd1 vccd1 _6036_/A sky130_fd_sc_hd__a21oi_2
XFILLER_98_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7986_ _7986_/A _8003_/B vssd1 vssd1 vccd1 vccd1 _7986_/X sky130_fd_sc_hd__or2_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9725_ _9893_/CLK _9725_/D vssd1 vssd1 vccd1 vccd1 _9725_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6937_ _6934_/X _6935_/X _6713_/C _6936_/X vssd1 vssd1 vccd1 vccd1 _6937_/X sky130_fd_sc_hd__o22a_1
XPHY_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9656_ _9656_/CLK _9656_/D vssd1 vssd1 vccd1 vccd1 _9656_/Q sky130_fd_sc_hd__dfxtp_1
X_6868_ _6868_/A _6868_/B vssd1 vssd1 vccd1 vccd1 _6868_/X sky130_fd_sc_hd__or2_1
X_8607_ _8574_/X _8577_/X _8561_/X _8578_/X vssd1 vssd1 vccd1 vccd1 _8623_/A sky130_fd_sc_hd__o22a_1
XFILLER_179_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9587_ _9923_/CLK _9587_/D vssd1 vssd1 vccd1 vccd1 _9587_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5819_ _5833_/A vssd1 vssd1 vccd1 vccd1 _5819_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8538_ _8610_/C _8538_/B vssd1 vssd1 vccd1 vccd1 _8573_/A sky130_fd_sc_hd__or2_1
X_6799_ _6797_/X _6798_/X _6797_/X _6798_/X vssd1 vssd1 vccd1 vccd1 _6806_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_157_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8469_ _8606_/A _8469_/B vssd1 vssd1 vccd1 vccd1 _8516_/A sky130_fd_sc_hd__or2_2
XFILLER_175_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7840_ _7840_/A _7840_/B vssd1 vssd1 vccd1 vccd1 _7844_/B sky130_fd_sc_hd__or2_1
X_7771_ _9927_/Q _6342_/Y _4802_/A _6350_/Y _7770_/X vssd1 vssd1 vccd1 vccd1 _7772_/D
+ sky130_fd_sc_hd__o221a_1
X_4983_ _5030_/A vssd1 vssd1 vccd1 vccd1 _5028_/A sky130_fd_sc_hd__inv_2
XFILLER_91_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6722_ _6722_/A vssd1 vssd1 vccd1 vccd1 _6723_/C sky130_fd_sc_hd__inv_2
X_9510_ _9527_/Q _9012_/X _7936_/Y _9014_/X _8970_/X _9053_/S vssd1 vssd1 vccd1 vccd1
+ _9510_/X sky130_fd_sc_hd__mux4_2
X_9441_ _9440_/X _6344_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _9441_/X sky130_fd_sc_hd__mux2_1
X_6653_ _6981_/A _6969_/B _6653_/C vssd1 vssd1 vccd1 vccd1 _6653_/X sky130_fd_sc_hd__or3_1
XFILLER_176_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5604_ _5604_/A vssd1 vssd1 vccd1 vccd1 _5604_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6584_ _6582_/X _6559_/Y _6576_/B vssd1 vssd1 vccd1 vccd1 _6584_/Y sky130_fd_sc_hd__o21ai_1
X_9372_ _7986_/X _6064_/Y _9504_/S vssd1 vssd1 vccd1 vccd1 _9372_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8323_ _4847_/X _8052_/Y _8373_/C _8322_/Y vssd1 vssd1 vccd1 vccd1 _8323_/X sky130_fd_sc_hd__o22a_1
X_5535_ _9476_/X _5489_/X _5587_/A vssd1 vssd1 vccd1 vccd1 _5582_/B sky130_fd_sc_hd__o21ai_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8254_ _9897_/Q _8254_/B vssd1 vssd1 vccd1 vccd1 _8254_/X sky130_fd_sc_hd__or2_1
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5466_ _9338_/X _9468_/X vssd1 vssd1 vccd1 vccd1 _5467_/B sky130_fd_sc_hd__nand2_1
XFILLER_132_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7205_ _7204_/A _7204_/B _7204_/X vssd1 vssd1 vccd1 vccd1 _7205_/X sky130_fd_sc_hd__a21bo_1
XFILLER_207_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8185_ _6365_/Y _9749_/Q _9845_/Q _7765_/Y vssd1 vssd1 vccd1 vccd1 _8187_/A sky130_fd_sc_hd__a22o_1
XFILLER_132_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5397_ _9716_/Q vssd1 vssd1 vccd1 vccd1 _5397_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7136_ _9424_/X vssd1 vssd1 vccd1 vccd1 _7169_/B sky130_fd_sc_hd__clkbuf_2
X_7067_ _6573_/X _6978_/A _7054_/B vssd1 vssd1 vccd1 vccd1 _7068_/A sky130_fd_sc_hd__o21ai_4
X_6018_ _6018_/A vssd1 vssd1 vccd1 vccd1 _6018_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7969_ _7969_/A _7981_/B vssd1 vssd1 vccd1 vccd1 _7969_/X sky130_fd_sc_hd__or2_1
XFILLER_14_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9708_ _9708_/CLK _9708_/D vssd1 vssd1 vccd1 vccd1 _9708_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9639_ _9828_/CLK _9639_/D vssd1 vssd1 vccd1 vccd1 _9639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5320_ _9724_/Q vssd1 vssd1 vccd1 vccd1 _5331_/A sky130_fd_sc_hd__inv_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5251_ _9746_/Q _5251_/B vssd1 vssd1 vccd1 vccd1 _5251_/Y sky130_fd_sc_hd__nand2_1
X_5182_ _5181_/X _5178_/X input26/X _5179_/X _5175_/X vssd1 vssd1 vccd1 vccd1 _9767_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8941_ _8938_/X _8940_/Y _8938_/X _8940_/Y vssd1 vssd1 vccd1 vccd1 _8941_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8872_ _8872_/A vssd1 vssd1 vccd1 vccd1 _8872_/Y sky130_fd_sc_hd__inv_2
X_7823_ _7823_/A _7823_/B vssd1 vssd1 vccd1 vccd1 _7827_/B sky130_fd_sc_hd__or2_1
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7754_ _7754_/A vssd1 vssd1 vccd1 vccd1 _7819_/A sky130_fd_sc_hd__buf_1
X_4966_ _5029_/A vssd1 vssd1 vccd1 vccd1 _4969_/A sky130_fd_sc_hd__inv_2
X_6705_ _6730_/A _6705_/B _6883_/A _6730_/B vssd1 vssd1 vccd1 vccd1 _6705_/X sky130_fd_sc_hd__or4_4
XPHY_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7685_ _8301_/A _7685_/B vssd1 vssd1 vccd1 vccd1 _9331_/S sky130_fd_sc_hd__nor2_2
X_4897_ _5631_/A vssd1 vssd1 vccd1 vccd1 _4897_/X sky130_fd_sc_hd__buf_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9424_ _7117_/X _5779_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9424_/X sky130_fd_sc_hd__mux2_2
X_6636_ _6807_/A vssd1 vssd1 vccd1 vccd1 _6760_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_192_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6567_ _6567_/A vssd1 vssd1 vccd1 vccd1 _6567_/Y sky130_fd_sc_hd__inv_2
X_9355_ _7064_/A _7622_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9355_/X sky130_fd_sc_hd__mux2_1
X_5518_ _5627_/A _8436_/C vssd1 vssd1 vccd1 vccd1 _5626_/A sky130_fd_sc_hd__or2_1
X_8306_ _9541_/Q vssd1 vssd1 vccd1 vccd1 _8306_/Y sky130_fd_sc_hd__inv_2
X_6498_ _6489_/X _6495_/X _6466_/Y _9796_/Q _6533_/B vssd1 vssd1 vccd1 vccd1 _6499_/A
+ sky130_fd_sc_hd__o32a_1
X_9286_ _9285_/X input23/X _9294_/S vssd1 vssd1 vccd1 vccd1 _9286_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8237_ _9755_/Q _8246_/A vssd1 vssd1 vccd1 vccd1 _8238_/B sky130_fd_sc_hd__or2_2
X_5449_ _6755_/A vssd1 vssd1 vccd1 vccd1 _6642_/A sky130_fd_sc_hd__clkbuf_2
X_8168_ _7680_/A _8097_/Y _9924_/Q _8096_/Y _8167_/X vssd1 vssd1 vccd1 vccd1 _8168_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_154_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7119_ _7107_/A _7107_/B _7108_/B vssd1 vssd1 vccd1 vccd1 _7119_/X sky130_fd_sc_hd__a21bo_1
XFILLER_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8099_ _9553_/Q _8081_/B _8082_/B vssd1 vssd1 vccd1 vccd1 _8099_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_47_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4820_ _7666_/A vssd1 vssd1 vccd1 vccd1 _4820_/X sky130_fd_sc_hd__buf_2
XFILLER_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4751_ _5918_/A _5147_/A _5844_/A vssd1 vssd1 vccd1 vccd1 _9282_/S sky130_fd_sc_hd__nor3_4
XFILLER_14_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7470_ _7470_/A _7470_/B vssd1 vssd1 vccd1 vccd1 _7470_/Y sky130_fd_sc_hd__nand2_2
XFILLER_174_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6421_ _6350_/A _8215_/A _6418_/Y vssd1 vssd1 vccd1 vccd1 _6538_/B sky130_fd_sc_hd__a21oi_2
XFILLER_119_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9140_ _9878_/Q _9894_/Q _9896_/Q vssd1 vssd1 vccd1 vccd1 _9140_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6352_ _9765_/Q vssd1 vssd1 vccd1 vccd1 _6352_/Y sky130_fd_sc_hd__inv_2
X_6283_ _9591_/Q vssd1 vssd1 vccd1 vccd1 _8040_/A sky130_fd_sc_hd__inv_2
X_9071_ _9070_/X _6349_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _9071_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5303_ _5299_/B _5224_/A _5302_/X _5275_/A _5240_/C vssd1 vssd1 vccd1 vccd1 _5304_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8022_ _9436_/X _8022_/B vssd1 vssd1 vccd1 vccd1 _8022_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5234_ _9736_/Q vssd1 vssd1 vccd1 vccd1 _5241_/A sky130_fd_sc_hd__inv_2
X_5165_ _5165_/A vssd1 vssd1 vccd1 vccd1 _5165_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5096_ _9833_/Q vssd1 vssd1 vccd1 vccd1 _5096_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8924_ _8922_/X _8923_/X _8922_/X _8923_/X vssd1 vssd1 vccd1 vccd1 _8924_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8855_ _8801_/A _8803_/Y _8804_/X _8808_/X vssd1 vssd1 vccd1 vccd1 _8895_/B sky130_fd_sc_hd__o22ai_2
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7806_ _4832_/X _7661_/B _7805_/Y vssd1 vssd1 vccd1 vccd1 _7806_/X sky130_fd_sc_hd__a21o_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8786_ _8787_/A _8787_/B vssd1 vssd1 vccd1 vccd1 _8786_/X sky130_fd_sc_hd__and2_1
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _5998_/A _5998_/B vssd1 vssd1 vccd1 vccd1 _5998_/X sky130_fd_sc_hd__or2_1
XFILLER_24_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7737_ _7852_/A vssd1 vssd1 vccd1 vccd1 _7738_/A sky130_fd_sc_hd__buf_1
XFILLER_24_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4949_ _9118_/X _4943_/X _9855_/Q _4944_/X _4947_/X vssd1 vssd1 vccd1 vccd1 _9855_/D
+ sky130_fd_sc_hd__o221a_1
X_7668_ _9911_/Q _7829_/A vssd1 vssd1 vccd1 vccd1 _7669_/B sky130_fd_sc_hd__or2_1
XFILLER_177_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6619_ _6969_/A _6660_/B vssd1 vssd1 vccd1 vccd1 _6620_/A sky130_fd_sc_hd__or2_2
X_9407_ _9406_/X _7005_/A _9507_/S vssd1 vssd1 vccd1 vccd1 _9407_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7599_ _7599_/A _7599_/B vssd1 vssd1 vccd1 vccd1 _7600_/B sky130_fd_sc_hd__or2_1
X_9338_ _7605_/Y _7560_/X _9475_/S vssd1 vssd1 vccd1 vccd1 _9338_/X sky130_fd_sc_hd__mux2_4
XFILLER_180_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9269_ _9268_/X _7825_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9269_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6970_ _6970_/A vssd1 vssd1 vccd1 vccd1 _6970_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5921_ _5937_/A vssd1 vssd1 vccd1 vccd1 _5921_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8640_ _8593_/Y _8596_/Y _8639_/X vssd1 vssd1 vccd1 vccd1 _8640_/Y sky130_fd_sc_hd__o21ai_2
X_5852_ _9631_/Q vssd1 vssd1 vccd1 vccd1 _5852_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8571_ _8571_/A _8571_/B vssd1 vssd1 vccd1 vccd1 _8619_/A sky130_fd_sc_hd__nor2_2
X_4803_ _9294_/X _4796_/X _4802_/X _4799_/X _4791_/X vssd1 vssd1 vccd1 vccd1 _9917_/D
+ sky130_fd_sc_hd__o221a_1
X_5783_ _9660_/Q _5774_/X _5769_/X _7108_/A _5772_/X vssd1 vssd1 vccd1 vccd1 _9660_/D
+ sky130_fd_sc_hd__o221a_1
X_7522_ _7522_/A _7522_/B vssd1 vssd1 vccd1 vccd1 _7522_/X sky130_fd_sc_hd__or2_1
XFILLER_21_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7453_ _7450_/X _7451_/X _7230_/C _7452_/X vssd1 vssd1 vccd1 vccd1 _7453_/X sky130_fd_sc_hd__o22a_1
X_6404_ _8200_/A _8199_/A _6402_/Y vssd1 vssd1 vccd1 vccd1 _6547_/B sky130_fd_sc_hd__a21oi_4
XFILLER_162_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7384_ _7384_/A _7384_/B _7384_/C _7407_/B vssd1 vssd1 vccd1 vccd1 _7384_/X sky130_fd_sc_hd__or4_4
XFILLER_115_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6335_ _6335_/A vssd1 vssd1 vccd1 vccd1 _6335_/Y sky130_fd_sc_hd__inv_2
X_9123_ _9607_/Q input19/X _9667_/Q vssd1 vssd1 vccd1 vccd1 _9123_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9054_ _8014_/Y _8013_/Y _9069_/S vssd1 vssd1 vccd1 vccd1 _9054_/X sky130_fd_sc_hd__mux2_1
X_6266_ _8027_/A _6140_/A _8029_/A _6245_/X _6256_/X vssd1 vssd1 vccd1 vccd1 _6266_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_130_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8005_ _8005_/A _8010_/B vssd1 vssd1 vccd1 vccd1 _8005_/Y sky130_fd_sc_hd__nor2_1
X_5217_ _4860_/X _5151_/X _8184_/B _5152_/X _5214_/X vssd1 vssd1 vccd1 vccd1 _9750_/D
+ sky130_fd_sc_hd__a221o_1
X_6197_ _6197_/A vssd1 vssd1 vccd1 vccd1 _6201_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5148_ _5882_/A _7922_/A vssd1 vssd1 vccd1 vccd1 _5179_/A sky130_fd_sc_hd__or2_4
XFILLER_84_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5079_ _5092_/A _5079_/B vssd1 vssd1 vccd1 vccd1 _9805_/D sky130_fd_sc_hd__nor2_1
XFILLER_151_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8907_ _8902_/X _8906_/Y _8902_/X _8906_/Y vssd1 vssd1 vccd1 vccd1 _8907_/X sky130_fd_sc_hd__a2bb2o_2
X_9887_ _9887_/CLK _9887_/D vssd1 vssd1 vccd1 vccd1 _9887_/Q sky130_fd_sc_hd__dfxtp_1
X_8838_ _8763_/X _8789_/X _8749_/X _8790_/X vssd1 vssd1 vccd1 vccd1 _8838_/X sky130_fd_sc_hd__o22a_1
X_8769_ _8708_/X _8709_/X _8703_/X _8707_/X vssd1 vssd1 vccd1 vccd1 _8769_/X sky130_fd_sc_hd__o211a_1
XFILLER_12_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6120_ _7121_/A vssd1 vssd1 vccd1 vccd1 _6120_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6051_ _6048_/A _6045_/X _6048_/A _6045_/X vssd1 vssd1 vccd1 vccd1 _6051_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5002_ _9834_/Q _4994_/X input30/X _4995_/X _5000_/X vssd1 vssd1 vccd1 vccd1 _9834_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9810_ _9928_/CLK _9810_/D vssd1 vssd1 vccd1 vccd1 _9810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9741_ _9887_/CLK _9741_/D vssd1 vssd1 vccd1 vccd1 _9741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6953_ _6943_/X _6944_/X _6945_/X _6952_/X vssd1 vssd1 vccd1 vccd1 _6954_/B sky130_fd_sc_hd__o22ai_2
XFILLER_207_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9672_ _9699_/CLK _9672_/D vssd1 vssd1 vccd1 vccd1 _9672_/Q sky130_fd_sc_hd__dfxtp_2
X_6884_ _6880_/X _6883_/X _6880_/X _6883_/X vssd1 vssd1 vccd1 vccd1 _6884_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5904_ _5910_/A vssd1 vssd1 vccd1 vccd1 _5909_/A sky130_fd_sc_hd__buf_1
X_8623_ _8623_/A _8623_/B vssd1 vssd1 vccd1 vccd1 _8709_/A sky130_fd_sc_hd__or2_1
X_5835_ _9641_/Q _5832_/X _5029_/X _5833_/X _5830_/X vssd1 vssd1 vccd1 vccd1 _9641_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8554_ _8554_/A vssd1 vssd1 vccd1 vccd1 _8555_/B sky130_fd_sc_hd__inv_2
X_5766_ _8381_/B _9664_/Q _5715_/Y vssd1 vssd1 vccd1 vccd1 _5766_/X sky130_fd_sc_hd__a21o_1
X_8485_ _8485_/A vssd1 vssd1 vccd1 vccd1 _8486_/B sky130_fd_sc_hd__inv_2
XFILLER_147_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5697_ _8967_/B vssd1 vssd1 vccd1 vccd1 _5697_/X sky130_fd_sc_hd__clkbuf_2
X_7505_ _7494_/A _7522_/B _7234_/A _7490_/B vssd1 vssd1 vccd1 vccd1 _7506_/B sky130_fd_sc_hd__o22a_1
XFILLER_107_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7436_ _7432_/X _7433_/X _7434_/X _7435_/X vssd1 vssd1 vccd1 vccd1 _7477_/B sky130_fd_sc_hd__o22a_1
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9106_ _6078_/X _6080_/X _9896_/Q vssd1 vssd1 vccd1 vccd1 _9106_/X sky130_fd_sc_hd__mux2_2
X_7367_ _7367_/A _7367_/B vssd1 vssd1 vccd1 vccd1 _7367_/X sky130_fd_sc_hd__or2_1
X_6318_ _6318_/A _6318_/B _6318_/C _6318_/D vssd1 vssd1 vccd1 vccd1 _6318_/X sky130_fd_sc_hd__and4_1
XFILLER_143_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7298_ _7298_/A _7304_/A vssd1 vssd1 vccd1 vccd1 _7298_/Y sky130_fd_sc_hd__nor2_1
X_6249_ _6265_/A _6248_/Y _6243_/A _6248_/A vssd1 vssd1 vccd1 vccd1 _6249_/X sky130_fd_sc_hd__o22a_1
X_9037_ _7987_/Y _9036_/X _9052_/S vssd1 vssd1 vccd1 vccd1 _9037_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5620_ _8176_/A _5620_/B vssd1 vssd1 vccd1 vccd1 _9702_/D sky130_fd_sc_hd__nor2_1
XFILLER_149_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5551_ _5549_/A _5548_/Y _9350_/S _5548_/A _5704_/A vssd1 vssd1 vccd1 vccd1 _5551_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_191_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8270_ _7819_/A _8242_/X _7726_/A _8244_/Y _8269_/X vssd1 vssd1 vccd1 vccd1 _8270_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_8_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5482_ _9394_/X _5481_/X _9394_/X _5481_/X vssd1 vssd1 vccd1 vccd1 _5482_/X sky130_fd_sc_hd__a2bb2o_1
X_7221_ _7359_/A vssd1 vssd1 vccd1 vccd1 _7247_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_6_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7152_ _7152_/A _7151_/X vssd1 vssd1 vccd1 vccd1 _7152_/X sky130_fd_sc_hd__or2b_1
XFILLER_140_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6103_ _6103_/A vssd1 vssd1 vccd1 vccd1 _6103_/X sky130_fd_sc_hd__buf_1
X_7083_ _7321_/D _7083_/B vssd1 vssd1 vccd1 vccd1 _7084_/B sky130_fd_sc_hd__or2_1
X_6034_ _9855_/Q _6034_/B vssd1 vssd1 vccd1 vccd1 _6034_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7985_ _8008_/B vssd1 vssd1 vccd1 vccd1 _8003_/B sky130_fd_sc_hd__buf_1
X_9724_ _9893_/CLK _9724_/D vssd1 vssd1 vccd1 vccd1 _9724_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6936_ _6934_/X _6935_/X _6934_/X _6935_/X vssd1 vssd1 vccd1 vccd1 _6936_/X sky130_fd_sc_hd__a2bb2o_1
XPHY_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9655_ _9656_/CLK _9655_/D vssd1 vssd1 vccd1 vccd1 _9655_/Q sky130_fd_sc_hd__dfxtp_1
X_6867_ _6867_/A _6867_/B _6867_/C _6867_/D vssd1 vssd1 vccd1 vccd1 _6867_/X sky130_fd_sc_hd__or4_4
XFILLER_194_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8606_ _8606_/A _8773_/B vssd1 vssd1 vccd1 vccd1 _8637_/A sky130_fd_sc_hd__or2_2
X_9586_ _9923_/CLK _9586_/D vssd1 vssd1 vccd1 vccd1 _9586_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5818_ _5832_/A vssd1 vssd1 vccd1 vccd1 _5818_/X sky130_fd_sc_hd__clkbuf_2
X_6798_ _6807_/A _9426_/X vssd1 vssd1 vccd1 vccd1 _6798_/X sky130_fd_sc_hd__or2_1
XFILLER_10_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8537_ _8535_/X _8536_/X _8535_/X _8536_/X vssd1 vssd1 vccd1 vccd1 _8538_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_194_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5749_ _9674_/Q _9657_/Q _5732_/Y _5748_/X vssd1 vssd1 vccd1 vccd1 _5749_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_22_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8468_ _8467_/A _8467_/B _8491_/A vssd1 vssd1 vccd1 vccd1 _8468_/X sky130_fd_sc_hd__a21bo_1
XFILLER_135_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8399_ _9686_/Q _6569_/Y _8432_/A _8398_/X vssd1 vssd1 vccd1 vccd1 _8399_/X sky130_fd_sc_hd__o22a_1
X_7419_ _7419_/A _7419_/B vssd1 vssd1 vccd1 vccd1 _7420_/B sky130_fd_sc_hd__or2_2
XFILLER_131_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput80 _9512_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_95_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7770_ _7865_/A _9769_/Q _7769_/Y _6341_/A vssd1 vssd1 vccd1 vccd1 _7770_/X sky130_fd_sc_hd__o22a_1
X_4982_ _5882_/A _9480_/S vssd1 vssd1 vccd1 vccd1 _5030_/A sky130_fd_sc_hd__or2_4
XFILLER_91_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6721_ _6730_/A _6721_/B vssd1 vssd1 vccd1 vccd1 _6722_/A sky130_fd_sc_hd__or2_2
X_9440_ _6316_/D _7897_/A _9480_/S vssd1 vssd1 vccd1 vccd1 _9440_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6652_ _6652_/A vssd1 vssd1 vccd1 vccd1 _6653_/C sky130_fd_sc_hd__inv_2
X_5603_ _5609_/A _5603_/B vssd1 vssd1 vccd1 vccd1 _9705_/D sky130_fd_sc_hd__nor2_1
X_9371_ _9370_/X _7005_/A _9507_/S vssd1 vssd1 vccd1 vccd1 _9371_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8322_ _8322_/A _9530_/Q vssd1 vssd1 vccd1 vccd1 _8322_/Y sky130_fd_sc_hd__nor2_1
X_6583_ _6576_/A _6576_/B _6577_/B vssd1 vssd1 vccd1 vccd1 _6583_/X sky130_fd_sc_hd__a21bo_1
X_5534_ _5588_/A _5588_/B vssd1 vssd1 vccd1 vccd1 _5587_/A sky130_fd_sc_hd__or2_1
XFILLER_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8253_ _8186_/A _9748_/Q _8187_/B vssd1 vssd1 vccd1 vccd1 _8254_/B sky130_fd_sc_hd__a21oi_1
X_5465_ _9338_/X _9468_/X vssd1 vssd1 vccd1 vccd1 _5467_/A sky130_fd_sc_hd__or2_1
X_8184_ _8184_/A _8184_/B vssd1 vssd1 vccd1 vccd1 _8184_/Y sky130_fd_sc_hd__nor2_1
XFILLER_132_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7204_ _7204_/A _7204_/B vssd1 vssd1 vccd1 vccd1 _7204_/X sky130_fd_sc_hd__or2_1
XFILLER_113_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7135_ _7490_/B vssd1 vssd1 vccd1 vccd1 _7135_/Y sky130_fd_sc_hd__inv_2
X_5396_ _9717_/Q vssd1 vssd1 vccd1 vccd1 _5396_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_clock/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7066_ _7066_/A vssd1 vssd1 vccd1 vccd1 _7071_/A sky130_fd_sc_hd__inv_2
XFILLER_100_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6017_ _6017_/A _6017_/B vssd1 vssd1 vccd1 vccd1 _6018_/A sky130_fd_sc_hd__or2_2
XFILLER_74_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7968_ _8773_/C vssd1 vssd1 vccd1 vccd1 _8955_/A sky130_fd_sc_hd__buf_6
XFILLER_14_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7899_ _7899_/A vssd1 vssd1 vccd1 vccd1 _7899_/Y sky130_fd_sc_hd__inv_2
XPHY_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9707_ _9828_/CLK _9707_/D vssd1 vssd1 vccd1 vccd1 _9707_/Q sky130_fd_sc_hd__dfxtp_1
X_6919_ _6915_/X _6916_/X _6917_/X _6918_/X vssd1 vssd1 vccd1 vccd1 _6919_/X sky130_fd_sc_hd__o22a_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9638_ _9650_/CLK _9638_/D vssd1 vssd1 vccd1 vccd1 _9638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9569_ _9888_/CLK _9569_/D vssd1 vssd1 vccd1 vccd1 _9569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5250_ _5250_/A _5259_/A vssd1 vssd1 vccd1 vccd1 _5251_/B sky130_fd_sc_hd__nor2_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5181_ _9767_/Q vssd1 vssd1 vccd1 vccd1 _5181_/X sky130_fd_sc_hd__buf_1
XFILLER_95_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8940_ _8940_/A vssd1 vssd1 vccd1 vccd1 _8940_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8871_ _8869_/Y _8904_/B _8869_/Y _8904_/B vssd1 vssd1 vccd1 vccd1 _8872_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7822_ _7665_/A _7665_/B _7821_/Y vssd1 vssd1 vccd1 vccd1 _7822_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7753_ _9907_/Q vssd1 vssd1 vccd1 vccd1 _7754_/A sky130_fd_sc_hd__inv_2
X_4965_ _4965_/A vssd1 vssd1 vccd1 vccd1 _9445_/S sky130_fd_sc_hd__inv_2
XFILLER_91_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6704_ _6842_/A vssd1 vssd1 vccd1 vccd1 _6730_/B sky130_fd_sc_hd__buf_1
XFILLER_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7684_ _7684_/A _7899_/A vssd1 vssd1 vccd1 vccd1 _7685_/B sky130_fd_sc_hd__or2_2
XFILLER_149_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9423_ _8966_/Y _8965_/Y _9490_/S vssd1 vssd1 vccd1 vccd1 _9423_/X sky130_fd_sc_hd__mux2_1
X_4896_ _5644_/A vssd1 vssd1 vccd1 vccd1 _5631_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_177_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6635_ _9612_/Q vssd1 vssd1 vccd1 vccd1 _6807_/A sky130_fd_sc_hd__inv_2
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6566_ _6564_/X _6565_/Y _6556_/B vssd1 vssd1 vccd1 vccd1 _6566_/Y sky130_fd_sc_hd__o21ai_1
X_9354_ _7633_/Y _7577_/X _9475_/S vssd1 vssd1 vccd1 vccd1 _9354_/X sky130_fd_sc_hd__mux2_2
X_5517_ _8452_/A _8416_/A vssd1 vssd1 vccd1 vccd1 _8436_/C sky130_fd_sc_hd__or2_2
XFILLER_180_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8305_ _9542_/Q vssd1 vssd1 vccd1 vccd1 _8305_/Y sky130_fd_sc_hd__inv_2
X_9285_ _9284_/X _7845_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9285_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8236_ _8236_/A _8236_/B vssd1 vssd1 vccd1 vccd1 _8246_/A sky130_fd_sc_hd__or2_1
X_6497_ _6500_/B vssd1 vssd1 vccd1 vccd1 _6533_/B sky130_fd_sc_hd__inv_2
XFILLER_105_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5448_ _6800_/A vssd1 vssd1 vccd1 vccd1 _6755_/A sky130_fd_sc_hd__clkbuf_2
X_8167_ _7680_/A _8097_/Y _4786_/X _8098_/Y _8166_/X vssd1 vssd1 vccd1 vccd1 _8167_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_120_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5379_ _5379_/A vssd1 vssd1 vccd1 vccd1 _5379_/X sky130_fd_sc_hd__clkbuf_2
X_8098_ _9554_/Q _8082_/B _8083_/B vssd1 vssd1 vccd1 vccd1 _8098_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_101_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7118_ _7108_/A _7108_/B _7109_/B vssd1 vssd1 vccd1 vccd1 _7118_/X sky130_fd_sc_hd__a21bo_1
X_7049_ _6951_/A _6951_/B _6951_/X vssd1 vssd1 vccd1 vccd1 _7066_/A sky130_fd_sc_hd__a21bo_1
XFILLER_101_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4750_ input7/X _5815_/B _5815_/D vssd1 vssd1 vccd1 vccd1 _5844_/A sky130_fd_sc_hd__or3_4
XFILLER_14_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6420_ _6420_/A vssd1 vssd1 vccd1 vccd1 _6539_/B sky130_fd_sc_hd__inv_2
XFILLER_162_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6351_ _6351_/A vssd1 vssd1 vccd1 vccd1 _6351_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5302_ _5240_/A _5305_/A _5240_/C vssd1 vssd1 vccd1 vccd1 _5302_/X sky130_fd_sc_hd__o21a_1
X_6282_ _6285_/A _6281_/X _6285_/A _6281_/X vssd1 vssd1 vccd1 vccd1 _6282_/X sky130_fd_sc_hd__a2bb2o_1
X_9070_ _6318_/C _7865_/A _9480_/S vssd1 vssd1 vccd1 vccd1 _9070_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8021_ _8021_/A _8021_/B vssd1 vssd1 vccd1 vccd1 _8021_/Y sky130_fd_sc_hd__nor2_1
X_5233_ _9737_/Q vssd1 vssd1 vccd1 vccd1 _5242_/A sky130_fd_sc_hd__inv_2
X_5164_ _9774_/Q vssd1 vssd1 vccd1 vccd1 _8205_/A sky130_fd_sc_hd__buf_2
XFILLER_96_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5095_ _9801_/Q vssd1 vssd1 vccd1 vccd1 _6318_/C sky130_fd_sc_hd__inv_2
XFILLER_110_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8923_ _8863_/X _8873_/X _8874_/X _8878_/X vssd1 vssd1 vccd1 vccd1 _8923_/X sky130_fd_sc_hd__o22a_1
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8854_ _8852_/X _8853_/X _8852_/X _8853_/X vssd1 vssd1 vccd1 vccd1 _8854_/Y sky130_fd_sc_hd__a2bb2oi_2
XFILLER_140_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7805_ _7805_/A vssd1 vssd1 vccd1 vccd1 _7805_/Y sky130_fd_sc_hd__inv_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8785_ _8710_/X _8718_/X _8719_/X _8727_/X vssd1 vssd1 vccd1 vccd1 _8787_/B sky130_fd_sc_hd__o22a_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5997_ _9851_/Q _5997_/B vssd1 vssd1 vccd1 vccd1 _5998_/B sky130_fd_sc_hd__nor2_1
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7736_ _9915_/Q vssd1 vssd1 vccd1 vccd1 _7852_/A sky130_fd_sc_hd__inv_2
X_4948_ _9119_/X _4943_/X _9856_/Q _4944_/X _4947_/X vssd1 vssd1 vccd1 vccd1 _9856_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_137_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7667_ _9910_/Q _7667_/B vssd1 vssd1 vccd1 vccd1 _7829_/A sky130_fd_sc_hd__or2_1
X_4879_ _4879_/A vssd1 vssd1 vccd1 vccd1 _4879_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_177_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6618_ _9463_/X vssd1 vssd1 vccd1 vccd1 _6971_/B sky130_fd_sc_hd__buf_1
X_9406_ _9405_/X _7490_/A _9506_/S vssd1 vssd1 vccd1 vccd1 _9406_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7598_ _7598_/A _7598_/B vssd1 vssd1 vccd1 vccd1 _7599_/B sky130_fd_sc_hd__or2_1
XFILLER_192_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6549_ _6550_/A _6549_/B vssd1 vssd1 vccd1 vccd1 _6549_/Y sky130_fd_sc_hd__nor2_1
XFILLER_118_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9337_ _7627_/X _7588_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9337_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9268_ _9759_/Q _9267_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9268_/X sky130_fd_sc_hd__mux2_1
X_9199_ _6543_/Y _9804_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9553_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8219_ _8219_/A _8219_/B vssd1 vssd1 vccd1 vccd1 _8219_/X sky130_fd_sc_hd__or2_1
XFILLER_121_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5920_ _5958_/A vssd1 vssd1 vccd1 vccd1 _5937_/A sky130_fd_sc_hd__buf_4
XFILLER_0_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5851_ _9632_/Q _5847_/X _5032_/X _5848_/X _5840_/X vssd1 vssd1 vccd1 vccd1 _9632_/D
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_2_0_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_clock/X
+ sky130_fd_sc_hd__clkbuf_1
X_8570_ _8568_/X _8613_/A _8568_/X _8613_/A vssd1 vssd1 vccd1 vccd1 _8571_/B sky130_fd_sc_hd__o2bb2a_1
X_4802_ _4802_/A vssd1 vssd1 vccd1 vccd1 _4802_/X sky130_fd_sc_hd__buf_1
X_5782_ _5782_/A vssd1 vssd1 vccd1 vccd1 _7108_/A sky130_fd_sc_hd__inv_2
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7521_ _7168_/X _7171_/X _7172_/X _7193_/X _7151_/X vssd1 vssd1 vccd1 vccd1 _7521_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_147_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7452_ _7450_/X _7451_/X _7450_/X _7451_/X vssd1 vssd1 vccd1 vccd1 _7452_/X sky130_fd_sc_hd__a2bb2o_1
X_6403_ _6343_/Y _6402_/Y _8197_/A vssd1 vssd1 vccd1 vccd1 _6405_/A sky130_fd_sc_hd__o21ai_1
XFILLER_174_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7383_ _9475_/X vssd1 vssd1 vccd1 vccd1 _7384_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_162_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6334_ _9792_/Q vssd1 vssd1 vccd1 vccd1 _6334_/Y sky130_fd_sc_hd__inv_2
X_9122_ _9606_/Q input18/X _9667_/Q vssd1 vssd1 vccd1 vccd1 _9122_/X sky130_fd_sc_hd__mux2_1
X_6265_ _6265_/A _6265_/B _6265_/C _6265_/D vssd1 vssd1 vccd1 vccd1 _6265_/X sky130_fd_sc_hd__or4_4
XFILLER_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9053_ _8011_/X _9052_/X _9053_/S vssd1 vssd1 vccd1 vccd1 _9053_/X sky130_fd_sc_hd__mux2_1
X_5216_ _9750_/Q vssd1 vssd1 vccd1 vccd1 _8184_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_142_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8004_ _9402_/X _8009_/B vssd1 vssd1 vccd1 vccd1 _8004_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6196_ _9575_/Q vssd1 vssd1 vccd1 vccd1 _7997_/A sky130_fd_sc_hd__inv_2
XFILLER_111_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5147_ _5147_/A _7918_/B vssd1 vssd1 vccd1 vccd1 _7922_/A sky130_fd_sc_hd__or2_4
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5078_ _5061_/X _6317_/C _5077_/Y _5073_/X vssd1 vssd1 vccd1 vccd1 _5079_/B sky130_fd_sc_hd__o22a_1
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8906_ _8906_/A vssd1 vssd1 vccd1 vccd1 _8906_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9886_ _9888_/CLK _9886_/D vssd1 vssd1 vccd1 vccd1 _9886_/Q sky130_fd_sc_hd__dfxtp_1
X_8837_ _8816_/X _8836_/X _8816_/X _8836_/X vssd1 vssd1 vccd1 vccd1 _8837_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8768_ _8768_/A vssd1 vssd1 vccd1 vccd1 _8893_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_157_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7719_ _9906_/Q _6339_/Y _9923_/Q _6345_/Y vssd1 vssd1 vccd1 vccd1 _7719_/X sky130_fd_sc_hd__o22a_1
XFILLER_8_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8699_ _8699_/A _8699_/B vssd1 vssd1 vccd1 vccd1 _8747_/A sky130_fd_sc_hd__nor2_2
XFILLER_165_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6050_ _6048_/A _6048_/B _6049_/Y vssd1 vssd1 vccd1 vccd1 _6050_/Y sky130_fd_sc_hd__a21oi_1
X_5001_ _9835_/Q _4994_/X input31/X _4995_/X _5000_/X vssd1 vssd1 vccd1 vccd1 _9835_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9740_ _9887_/CLK _9740_/D vssd1 vssd1 vccd1 vccd1 _9740_/Q sky130_fd_sc_hd__dfxtp_1
X_6952_ _6946_/X _6948_/X _6949_/X _6951_/X vssd1 vssd1 vccd1 vccd1 _6952_/X sky130_fd_sc_hd__o22a_1
XFILLER_201_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9671_ _9673_/CLK _9671_/D vssd1 vssd1 vccd1 vccd1 _9671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6883_ _6883_/A _6883_/B _6883_/C vssd1 vssd1 vccd1 vccd1 _6883_/X sky130_fd_sc_hd__or3_1
X_5903_ _5903_/A _9138_/X vssd1 vssd1 vccd1 vccd1 _9606_/D sky130_fd_sc_hd__and2_1
X_8622_ _8621_/A _8620_/Y _8621_/Y _8620_/A vssd1 vssd1 vccd1 vccd1 _8623_/B sky130_fd_sc_hd__a22o_1
X_5834_ _9642_/Q _5832_/X _5026_/X _5833_/X _5830_/X vssd1 vssd1 vccd1 vccd1 _9642_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8553_ _8551_/X _8552_/X _8551_/X _8552_/X vssd1 vssd1 vccd1 vccd1 _8554_/A sky130_fd_sc_hd__a2bb2o_2
X_5765_ _9665_/Q _5697_/X _5570_/X _5764_/Y _5698_/X vssd1 vssd1 vccd1 vccd1 _9665_/D
+ sky130_fd_sc_hd__o221a_1
X_8484_ _8516_/A _8483_/B _8483_/X vssd1 vssd1 vccd1 vccd1 _8485_/A sky130_fd_sc_hd__a21bo_1
XFILLER_147_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5696_ _6569_/A _5689_/X _9097_/X _5692_/X _5690_/X vssd1 vssd1 vccd1 vccd1 _9670_/D
+ sky130_fd_sc_hd__o221a_1
X_7504_ _7501_/X _7503_/X _7501_/X _7503_/X vssd1 vssd1 vccd1 vccd1 _7504_/X sky130_fd_sc_hd__a2bb2o_1
X_7435_ _7432_/X _7433_/X _7432_/X _7433_/X vssd1 vssd1 vccd1 vccd1 _7435_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7366_ _7348_/B _7350_/B _7348_/B _7365_/X vssd1 vssd1 vccd1 vccd1 _7367_/B sky130_fd_sc_hd__a2bb2o_1
X_6317_ _6317_/A _6317_/B _6317_/C _6317_/D vssd1 vssd1 vccd1 vccd1 _6317_/X sky130_fd_sc_hd__and4_1
X_9105_ _6069_/X _6072_/X _9896_/Q vssd1 vssd1 vccd1 vccd1 _9105_/X sky130_fd_sc_hd__mux2_2
XFILLER_1_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7297_ _7282_/A _7292_/Y _7289_/X _7293_/X vssd1 vssd1 vccd1 vccd1 _7304_/A sky130_fd_sc_hd__o22ai_4
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6248_ _6248_/A vssd1 vssd1 vccd1 vccd1 _6248_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9036_ _7988_/Y _9605_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9036_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6179_ _6179_/A _6179_/B vssd1 vssd1 vccd1 vccd1 _6187_/A sky130_fd_sc_hd__or2_1
XFILLER_97_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9869_ _9895_/CLK _9869_/D vssd1 vssd1 vccd1 vccd1 _9869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5550_ _5586_/A vssd1 vssd1 vccd1 vccd1 _5704_/A sky130_fd_sc_hd__buf_2
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5481_ _5479_/Y _5480_/Y _5479_/Y _5480_/Y vssd1 vssd1 vccd1 vccd1 _5481_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_8_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7220_ _9472_/X vssd1 vssd1 vccd1 vccd1 _7359_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_144_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7151_ _7178_/A _7494_/B _7491_/A _7169_/B vssd1 vssd1 vccd1 vccd1 _7151_/X sky130_fd_sc_hd__or4_4
XFILLER_98_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7082_ _7038_/Y _7081_/X _7038_/Y _7081_/X vssd1 vssd1 vccd1 vccd1 _7082_/Y sky130_fd_sc_hd__a2bb2oi_1
X_6102_ _8003_/A _9649_/Q _9862_/Q _6101_/Y vssd1 vssd1 vccd1 vccd1 _6103_/A sky130_fd_sc_hd__a22o_1
XFILLER_140_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6033_ _9642_/Q vssd1 vssd1 vccd1 vccd1 _6034_/B sky130_fd_sc_hd__inv_2
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7984_ _9367_/X _8002_/B vssd1 vssd1 vccd1 vccd1 _7984_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9723_ _9893_/CLK _9723_/D vssd1 vssd1 vccd1 vccd1 _9723_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6935_ _6926_/A _6926_/B _6926_/X vssd1 vssd1 vccd1 vccd1 _6935_/X sky130_fd_sc_hd__a21bo_1
XFILLER_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6866_ _9427_/X vssd1 vssd1 vccd1 vccd1 _6867_/B sky130_fd_sc_hd__buf_2
X_9654_ _9673_/CLK _9654_/D vssd1 vssd1 vccd1 vccd1 _9654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9585_ _9836_/CLK _9585_/D vssd1 vssd1 vccd1 vccd1 _9585_/Q sky130_fd_sc_hd__dfxtp_1
X_8605_ _8605_/A _9392_/X vssd1 vssd1 vccd1 vccd1 _8686_/A sky130_fd_sc_hd__or2_2
XPHY_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5817_ _5833_/A vssd1 vssd1 vccd1 vccd1 _5832_/A sky130_fd_sc_hd__inv_2
X_6797_ _6800_/A _9425_/X vssd1 vssd1 vccd1 vccd1 _6797_/X sky130_fd_sc_hd__or2_1
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8536_ _8566_/A _9382_/X _8536_/C vssd1 vssd1 vccd1 vccd1 _8536_/X sky130_fd_sc_hd__or3_1
XFILLER_194_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5748_ _8391_/B _5735_/Y _5736_/X _5747_/X vssd1 vssd1 vccd1 vccd1 _5748_/X sky130_fd_sc_hd__o22a_1
XFILLER_10_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8467_ _8467_/A _8467_/B vssd1 vssd1 vccd1 vccd1 _8491_/A sky130_fd_sc_hd__or2_1
XFILLER_135_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5679_ _6593_/A _5671_/X _9108_/X _5676_/X _5674_/X vssd1 vssd1 vccd1 vccd1 _9681_/D
+ sky130_fd_sc_hd__o221a_1
X_8398_ _9685_/Q _6571_/Y _8397_/Y vssd1 vssd1 vccd1 vccd1 _8398_/X sky130_fd_sc_hd__o21ba_1
X_7418_ _7394_/C _7391_/B _7391_/Y vssd1 vssd1 vccd1 vccd1 _7419_/B sky130_fd_sc_hd__o21ai_1
XFILLER_190_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7349_ _7337_/X _7338_/X _7337_/X _7338_/X vssd1 vssd1 vccd1 vccd1 _7350_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_173_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9019_ _9018_/X _9752_/Q _9481_/S vssd1 vssd1 vccd1 vccd1 _9019_/X sky130_fd_sc_hd__mux2_2
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput70 _9062_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_110_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput81 _9513_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4981_ _5815_/A _5815_/B _9038_/S vssd1 vssd1 vccd1 vccd1 _9480_/S sky130_fd_sc_hd__or3_4
XFILLER_51_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6720_ _6701_/X _6705_/X _6718_/X _6719_/X vssd1 vssd1 vccd1 vccd1 _6720_/X sky130_fd_sc_hd__o22a_1
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6651_ _6975_/A _7006_/B vssd1 vssd1 vccd1 vccd1 _6652_/A sky130_fd_sc_hd__or2_2
X_5602_ _5586_/X _5599_/Y _5600_/Y _7642_/A _5577_/X vssd1 vssd1 vccd1 vccd1 _5603_/B
+ sky130_fd_sc_hd__o32a_1
X_6582_ _6582_/A vssd1 vssd1 vccd1 vccd1 _6582_/X sky130_fd_sc_hd__clkbuf_2
X_9370_ _9369_/X _7490_/A _9506_/S vssd1 vssd1 vccd1 vccd1 _9370_/X sky130_fd_sc_hd__mux2_1
X_8321_ _8322_/A _9530_/Q _7778_/B _9529_/Q vssd1 vssd1 vccd1 vccd1 _8373_/C sky130_fd_sc_hd__a22oi_2
X_5533_ _9428_/X _5493_/X _5494_/X _5532_/X vssd1 vssd1 vccd1 vccd1 _5588_/B sky130_fd_sc_hd__o22a_1
XFILLER_117_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8252_ _8188_/Y _8251_/X _8188_/Y _8251_/X vssd1 vssd1 vccd1 vccd1 _8252_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_117_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5464_ _9340_/X _9339_/X _5406_/X _5463_/X vssd1 vssd1 vccd1 vccd1 _5464_/Y sky130_fd_sc_hd__o22ai_1
X_8183_ _8183_/A _8183_/B vssd1 vssd1 vccd1 vccd1 _8183_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7203_ _7518_/A _9432_/X _7202_/X vssd1 vssd1 vccd1 vccd1 _7204_/B sky130_fd_sc_hd__or3b_1
X_5395_ _5395_/A vssd1 vssd1 vccd1 vccd1 _9719_/D sky130_fd_sc_hd__inv_2
X_7134_ _7178_/B vssd1 vssd1 vccd1 vccd1 _7490_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_101_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7065_ _7065_/A vssd1 vssd1 vccd1 vccd1 _7072_/A sky130_fd_sc_hd__inv_2
XFILLER_100_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6016_ _7955_/A _9640_/Q vssd1 vssd1 vccd1 vccd1 _6017_/B sky130_fd_sc_hd__nor2_1
XFILLER_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7967_ _7967_/A vssd1 vssd1 vccd1 vccd1 _8773_/C sky130_fd_sc_hd__clkbuf_2
XPHY_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7898_ _4775_/X _7893_/Y _7860_/X _7902_/B vssd1 vssd1 vccd1 vccd1 _7898_/X sky130_fd_sc_hd__o211a_1
XPHY_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9706_ _9708_/CLK _9706_/D vssd1 vssd1 vccd1 vccd1 _9706_/Q sky130_fd_sc_hd__dfxtp_1
X_6918_ _6915_/X _6916_/X _6915_/X _6916_/X vssd1 vssd1 vccd1 vccd1 _6918_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_195_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9637_ _9828_/CLK _9637_/D vssd1 vssd1 vccd1 vccd1 _9637_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6849_ _6844_/X _6848_/X _6844_/X _6848_/X vssd1 vssd1 vccd1 vccd1 _6849_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_210_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9568_ _9888_/CLK _9568_/D vssd1 vssd1 vccd1 vccd1 _9568_/Q sky130_fd_sc_hd__dfxtp_1
X_8519_ _8515_/X _8518_/X _8515_/X _8518_/X vssd1 vssd1 vccd1 vccd1 _8519_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_108_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9499_ _7955_/X _6014_/B _9504_/S vssd1 vssd1 vccd1 vccd1 _9499_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5180_ _6350_/A _5178_/X input28/X _5179_/X _5175_/X vssd1 vssd1 vccd1 vccd1 _9768_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8870_ _8865_/C _8824_/Y _8825_/X _8830_/X vssd1 vssd1 vccd1 vccd1 _8904_/B sky130_fd_sc_hd__o22ai_2
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7821_ _7821_/A vssd1 vssd1 vccd1 vccd1 _7821_/Y sky130_fd_sc_hd__inv_2
X_7752_ _7752_/A _7752_/B _7752_/C _7752_/D vssd1 vssd1 vccd1 vccd1 _7773_/C sky130_fd_sc_hd__and4_1
X_4964_ _5816_/A _8047_/B vssd1 vssd1 vccd1 vccd1 _4965_/A sky130_fd_sc_hd__or2_2
XFILLER_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6703_ _9095_/X vssd1 vssd1 vccd1 vccd1 _6842_/A sky130_fd_sc_hd__clkbuf_2
X_7683_ _7683_/A _7683_/B vssd1 vssd1 vccd1 vccd1 _7899_/A sky130_fd_sc_hd__or2_1
X_9422_ _8846_/Y _8845_/B _9477_/S vssd1 vssd1 vccd1 vccd1 _9422_/X sky130_fd_sc_hd__mux2_2
X_4895_ _5348_/B vssd1 vssd1 vccd1 vccd1 _5644_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_177_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6634_ _6678_/A _9461_/X vssd1 vssd1 vccd1 vccd1 _6634_/X sky130_fd_sc_hd__or2_1
XFILLER_22_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6565_ _6565_/A vssd1 vssd1 vccd1 vccd1 _6565_/Y sky130_fd_sc_hd__inv_2
X_9353_ _7617_/X _7583_/A _9475_/S vssd1 vssd1 vccd1 vccd1 _9353_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6496_ _6353_/A _8225_/A _8223_/A vssd1 vssd1 vccd1 vccd1 _6500_/B sky130_fd_sc_hd__a21bo_1
X_5516_ _5515_/X _5442_/A _9684_/Q _5442_/A vssd1 vssd1 vccd1 vccd1 _8416_/A sky130_fd_sc_hd__o2bb2a_2
X_8304_ _4812_/X _8303_/Y _4814_/X _8111_/Y vssd1 vssd1 vccd1 vccd1 _8328_/A sky130_fd_sc_hd__a22o_1
X_9284_ _9764_/Q _9283_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9284_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8235_ _9753_/Q _8235_/B vssd1 vssd1 vccd1 vccd1 _8236_/B sky130_fd_sc_hd__or2_2
X_5447_ _9611_/Q vssd1 vssd1 vccd1 vccd1 _6800_/A sky130_fd_sc_hd__inv_2
XFILLER_160_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8166_ _4788_/X _8099_/Y _4786_/X _8098_/Y _8165_/X vssd1 vssd1 vccd1 vccd1 _8166_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5378_ _5378_/A vssd1 vssd1 vccd1 vccd1 _9723_/D sky130_fd_sc_hd__inv_2
XFILLER_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8097_ _9555_/Q _8083_/B _8084_/B vssd1 vssd1 vccd1 vccd1 _8097_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_120_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7117_ _7109_/A _7109_/B _7110_/B vssd1 vssd1 vccd1 vccd1 _7117_/X sky130_fd_sc_hd__a21bo_1
XFILLER_170_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7048_ _6949_/X _6951_/X _6949_/X _6951_/X vssd1 vssd1 vccd1 vccd1 _7065_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8999_ _9523_/Q _5041_/A _8999_/S vssd1 vssd1 vccd1 vccd1 _8999_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6350_ _6350_/A vssd1 vssd1 vccd1 vccd1 _6350_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5301_ _5301_/A vssd1 vssd1 vccd1 vccd1 _9736_/D sky130_fd_sc_hd__inv_2
X_6281_ _9589_/Q _6171_/A _6275_/X _6277_/Y vssd1 vssd1 vccd1 vccd1 _6281_/X sky130_fd_sc_hd__a22o_1
XFILLER_142_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8020_ _9391_/X _8030_/B vssd1 vssd1 vccd1 vccd1 _8020_/X sky130_fd_sc_hd__and2_1
XFILLER_115_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5232_ _9738_/Q vssd1 vssd1 vccd1 vccd1 _5243_/A sky130_fd_sc_hd__inv_2
X_5163_ _5162_/X _5155_/X input35/X _5157_/X _5153_/X vssd1 vssd1 vccd1 vccd1 _9775_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5094_ _8177_/A vssd1 vssd1 vccd1 vccd1 _5115_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_96_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8922_ _8915_/X _8921_/X _8915_/X _8921_/X vssd1 vssd1 vccd1 vccd1 _8922_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8853_ _8722_/A _8806_/A _8807_/A _8893_/B vssd1 vssd1 vccd1 vccd1 _8853_/X sky130_fd_sc_hd__a211o_2
X_7804_ _4835_/X _7798_/Y _7807_/B _7785_/X vssd1 vssd1 vccd1 vccd1 _7804_/X sky130_fd_sc_hd__o211a_1
XFILLER_169_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8784_ _8771_/X _8783_/X _8771_/X _8783_/X vssd1 vssd1 vccd1 vccd1 _8787_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _9638_/Q vssd1 vssd1 vccd1 vccd1 _5997_/B sky130_fd_sc_hd__inv_2
XFILLER_12_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7735_ _9925_/Q vssd1 vssd1 vccd1 vccd1 _7895_/A sky130_fd_sc_hd__inv_2
XFILLER_24_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4947_ _4991_/A vssd1 vssd1 vccd1 vccd1 _4947_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7666_ _7666_/A _7821_/A vssd1 vssd1 vccd1 vccd1 _7667_/B sky130_fd_sc_hd__or2_1
X_4878_ _9741_/Q _4870_/X _9889_/Q _4871_/X _4873_/X vssd1 vssd1 vccd1 vccd1 _9889_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_137_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6617_ _6707_/A vssd1 vssd1 vccd1 vccd1 _7006_/A sky130_fd_sc_hd__buf_2
X_9405_ _9404_/X _8955_/A _9505_/S vssd1 vssd1 vccd1 vccd1 _9405_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7597_ _7597_/A _7597_/B vssd1 vssd1 vccd1 vccd1 _7598_/B sky130_fd_sc_hd__or2_1
X_9336_ _7066_/A _7626_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9336_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6548_ _6550_/A _6548_/B vssd1 vssd1 vccd1 vccd1 _6548_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6479_ _9786_/Q _6520_/B _9785_/Q _6519_/B vssd1 vssd1 vccd1 vccd1 _6480_/B sky130_fd_sc_hd__o22ai_1
XFILLER_106_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9267_ _7822_/X _9759_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9267_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9198_ _6541_/Y _9803_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9552_/D sky130_fd_sc_hd__mux2_1
X_8218_ _6350_/A _8216_/B _8216_/Y vssd1 vssd1 vccd1 vccd1 _8218_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_133_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8149_ _7761_/X _8115_/X _8148_/X vssd1 vssd1 vccd1 vccd1 _8149_/Y sky130_fd_sc_hd__a21oi_1
XINSDIODE2_0 _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5850_ _9633_/Q _5847_/X _5029_/X _5848_/X _5840_/X vssd1 vssd1 vccd1 vccd1 _9633_/D
+ sky130_fd_sc_hd__o221a_1
X_4801_ _9917_/Q vssd1 vssd1 vccd1 vccd1 _4802_/A sky130_fd_sc_hd__clkbuf_2
X_5781_ _5727_/X _5751_/X _5727_/X _5751_/X vssd1 vssd1 vccd1 vccd1 _5782_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7520_ _7497_/X _7519_/Y _7497_/X _7519_/Y vssd1 vssd1 vccd1 vccd1 _7520_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_202_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7451_ _7443_/A _7443_/B _7443_/X vssd1 vssd1 vccd1 vccd1 _7451_/X sky130_fd_sc_hd__a21bo_1
X_6402_ _6402_/A vssd1 vssd1 vccd1 vccd1 _6402_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7382_ _7382_/A _7381_/X vssd1 vssd1 vccd1 vccd1 _7382_/X sky130_fd_sc_hd__or2b_1
X_6333_ _9761_/Q vssd1 vssd1 vccd1 vccd1 _6333_/Y sky130_fd_sc_hd__inv_2
X_9121_ _9605_/Q input17/X _9667_/Q vssd1 vssd1 vccd1 vccd1 _9121_/X sky130_fd_sc_hd__mux2_1
X_6264_ _9587_/Q _6170_/A _8031_/A _6140_/A vssd1 vssd1 vccd1 vccd1 _6268_/A sky130_fd_sc_hd__a22o_1
XFILLER_115_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9052_ _8009_/Y _9051_/X _9052_/S vssd1 vssd1 vccd1 vccd1 _9052_/X sky130_fd_sc_hd__mux2_2
X_5215_ _5035_/X _5151_/X _8183_/B _5152_/X _5214_/X vssd1 vssd1 vccd1 vccd1 _9751_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8003_ _8003_/A _8003_/B vssd1 vssd1 vccd1 vccd1 _8003_/X sky130_fd_sc_hd__or2_1
X_6195_ _6200_/B _6194_/Y _6200_/B _6194_/Y vssd1 vssd1 vccd1 vccd1 _6195_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5146_ _5815_/A input8/X _5815_/D vssd1 vssd1 vccd1 vccd1 _7918_/B sky130_fd_sc_hd__or3_4
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5077_ _9837_/Q vssd1 vssd1 vccd1 vccd1 _5077_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8905_ _8832_/A _8903_/Y _8872_/Y _8869_/Y _8904_/X vssd1 vssd1 vccd1 vccd1 _8906_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9885_ _9888_/CLK _9885_/D vssd1 vssd1 vccd1 vccd1 _9885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8836_ _8818_/X _8835_/X _8818_/X _8835_/X vssd1 vssd1 vccd1 vccd1 _8836_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8767_ _8711_/X _8712_/X _8713_/X _8717_/Y _8766_/X vssd1 vssd1 vccd1 vccd1 _8767_/X
+ sky130_fd_sc_hd__o221a_1
X_5979_ _9636_/Q vssd1 vssd1 vccd1 vccd1 _5979_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7718_ _9923_/Q vssd1 vssd1 vccd1 vccd1 _7887_/A sky130_fd_sc_hd__inv_2
XFILLER_40_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8698_ _8698_/A vssd1 vssd1 vccd1 vccd1 _8699_/B sky130_fd_sc_hd__inv_2
XFILLER_193_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7649_ _7652_/B _9711_/Q vssd1 vssd1 vccd1 vccd1 _7649_/Y sky130_fd_sc_hd__nor2b_1
XFILLER_20_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9319_ _7896_/Y _9776_/Q _9327_/S vssd1 vssd1 vccd1 vccd1 _9319_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5000_ _5036_/A vssd1 vssd1 vccd1 vccd1 _5000_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6951_ _6951_/A _6951_/B vssd1 vssd1 vccd1 vccd1 _6951_/X sky130_fd_sc_hd__or2_1
XFILLER_207_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9670_ _9673_/CLK _9670_/D vssd1 vssd1 vccd1 vccd1 _9670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5902_ _5903_/A _9072_/X vssd1 vssd1 vccd1 vccd1 _9607_/D sky130_fd_sc_hd__and2_1
X_6882_ _6882_/A vssd1 vssd1 vccd1 vccd1 _6883_/C sky130_fd_sc_hd__inv_2
X_8621_ _8621_/A vssd1 vssd1 vccd1 vccd1 _8621_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5833_ _5833_/A vssd1 vssd1 vccd1 vccd1 _5833_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8552_ _8515_/X _8518_/X _8483_/X _8519_/X vssd1 vssd1 vccd1 vccd1 _8552_/X sky130_fd_sc_hd__o22a_1
XFILLER_61_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5764_ _7492_/B vssd1 vssd1 vccd1 vccd1 _5764_/Y sky130_fd_sc_hd__inv_2
X_7503_ _7503_/A _7503_/B vssd1 vssd1 vccd1 vccd1 _7503_/X sky130_fd_sc_hd__or2_1
X_8483_ _8516_/A _8483_/B vssd1 vssd1 vccd1 vccd1 _8483_/X sky130_fd_sc_hd__or2_1
X_5695_ _8394_/B _5689_/X _9098_/X _5692_/X _5690_/X vssd1 vssd1 vccd1 vccd1 _9671_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_162_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7434_ _7259_/A _7259_/B _7260_/B vssd1 vssd1 vccd1 vccd1 _7434_/X sky130_fd_sc_hd__a21bo_1
XFILLER_162_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7365_ _7350_/A _7350_/B _7350_/X vssd1 vssd1 vccd1 vccd1 _7365_/X sky130_fd_sc_hd__a21bo_1
X_6316_ _6316_/A _6316_/B _6316_/C _6316_/D vssd1 vssd1 vccd1 vccd1 _6316_/X sky130_fd_sc_hd__and4_1
XFILLER_131_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9104_ _6060_/X _6062_/X _9896_/Q vssd1 vssd1 vccd1 vccd1 _9104_/X sky130_fd_sc_hd__mux2_2
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7296_ _7296_/A vssd1 vssd1 vccd1 vccd1 _7298_/A sky130_fd_sc_hd__inv_2
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6247_ _6247_/A _6247_/B vssd1 vssd1 vccd1 vccd1 _6248_/A sky130_fd_sc_hd__nand2_1
X_9035_ _7984_/Y _9034_/X _9038_/S vssd1 vssd1 vccd1 vccd1 _9035_/X sky130_fd_sc_hd__mux2_2
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6178_ _6152_/X _6155_/X _6176_/X _6160_/X _6177_/X vssd1 vssd1 vccd1 vccd1 _6179_/B
+ sky130_fd_sc_hd__o311a_1
X_5129_ _5128_/X _9791_/Q _5121_/X _9218_/X _5124_/X vssd1 vssd1 vccd1 vccd1 _9791_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9868_ _9874_/CLK _9868_/D vssd1 vssd1 vccd1 vccd1 _9868_/Q sky130_fd_sc_hd__dfxtp_1
X_8819_ _9429_/X vssd1 vssd1 vccd1 vccd1 _8942_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_111_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9799_ _9916_/CLK _9799_/D vssd1 vssd1 vccd1 vccd1 _9799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5480_ _5415_/A _5415_/B _5415_/Y vssd1 vssd1 vccd1 vccd1 _5480_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7150_ _7178_/A _7494_/B _7265_/A _7169_/B vssd1 vssd1 vccd1 vccd1 _7152_/A sky130_fd_sc_hd__o22a_1
X_7081_ _7081_/A _7081_/B vssd1 vssd1 vccd1 vccd1 _7081_/X sky130_fd_sc_hd__or2_1
X_6101_ _9649_/Q vssd1 vssd1 vccd1 vccd1 _6101_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6032_ _6026_/Y _6031_/A _6026_/A _6031_/Y vssd1 vssd1 vccd1 vccd1 _6032_/X sky130_fd_sc_hd__o22a_1
XFILLER_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7983_ _7983_/A _7993_/B vssd1 vssd1 vccd1 vccd1 _7983_/Y sky130_fd_sc_hd__nor2_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_9722_ _9893_/CLK _9722_/D vssd1 vssd1 vccd1 vccd1 _9722_/Q sky130_fd_sc_hd__dfxtp_1
X_6934_ _6857_/A _6857_/B _6859_/A vssd1 vssd1 vccd1 vccd1 _6934_/X sky130_fd_sc_hd__a21bo_1
XPHY_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9653_ _9673_/CLK _9653_/D vssd1 vssd1 vccd1 vccd1 _9653_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8604_ _8603_/A _8603_/B _8650_/A vssd1 vssd1 vccd1 vccd1 _8604_/X sky130_fd_sc_hd__a21bo_1
XPHY_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6865_ _6865_/A _6864_/X vssd1 vssd1 vccd1 vccd1 _6865_/X sky130_fd_sc_hd__or2b_1
XFILLER_194_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9584_ _9833_/CLK _9584_/D vssd1 vssd1 vccd1 vccd1 _9584_/Q sky130_fd_sc_hd__dfxtp_1
X_5816_ _5816_/A _7911_/A vssd1 vssd1 vccd1 vccd1 _5833_/A sky130_fd_sc_hd__or2_2
X_6796_ _6821_/B _9427_/X _6796_/C _6796_/D vssd1 vssd1 vccd1 vccd1 _6796_/X sky130_fd_sc_hd__or4_4
XFILLER_22_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8535_ _8605_/A _9457_/X vssd1 vssd1 vccd1 vccd1 _8535_/X sky130_fd_sc_hd__or2_2
X_5747_ _6564_/A _5738_/Y _5739_/X _5746_/X vssd1 vssd1 vccd1 vccd1 _5747_/X sky130_fd_sc_hd__o22a_1
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8466_ _8466_/A vssd1 vssd1 vccd1 vccd1 _8467_/B sky130_fd_sc_hd__inv_2
X_5678_ _6982_/A _5671_/X _9109_/X _5676_/X _5674_/X vssd1 vssd1 vccd1 vccd1 _9682_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_108_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7417_ _7405_/A _7405_/B _7442_/A vssd1 vssd1 vccd1 vccd1 _7420_/A sky130_fd_sc_hd__a21o_1
XFILLER_163_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8397_ _5515_/X _6890_/A _8396_/X vssd1 vssd1 vccd1 vccd1 _8397_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7348_ _7352_/B _7348_/B vssd1 vssd1 vccd1 vccd1 _7348_/X sky130_fd_sc_hd__and2b_1
XFILLER_131_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7279_ _7266_/Y _7267_/X _7266_/Y _7267_/X vssd1 vssd1 vccd1 vccd1 _7279_/X sky130_fd_sc_hd__a2bb2o_1
X_9018_ _9784_/Q _9901_/Q _9480_/S vssd1 vssd1 vccd1 vccd1 _9018_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput60 _9053_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[15] sky130_fd_sc_hd__clkbuf_2
Xoutput71 _9063_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput82 _9514_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4980_ _5918_/A vssd1 vssd1 vccd1 vccd1 _5882_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6650_ _6631_/X _6632_/X _6648_/X _6649_/X vssd1 vssd1 vccd1 vccd1 _6650_/X sky130_fd_sc_hd__o22a_1
X_5601_ _9705_/Q vssd1 vssd1 vccd1 vccd1 _7642_/A sky130_fd_sc_hd__inv_2
X_6581_ _6577_/A _6577_/B _6578_/B vssd1 vssd1 vccd1 vccd1 _6581_/X sky130_fd_sc_hd__a21bo_1
X_8320_ _8369_/A vssd1 vssd1 vccd1 vccd1 _8320_/Y sky130_fd_sc_hd__inv_2
X_5532_ _9403_/X _5497_/X _5594_/A vssd1 vssd1 vccd1 vccd1 _5532_/X sky130_fd_sc_hd__o21a_1
XFILLER_117_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8251_ _8184_/A _8184_/B _8184_/Y vssd1 vssd1 vccd1 vccd1 _8251_/X sky130_fd_sc_hd__a21o_1
XFILLER_145_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5463_ _9344_/X _9342_/X _5409_/Y _5471_/A vssd1 vssd1 vccd1 vccd1 _5463_/X sky130_fd_sc_hd__o22a_1
XFILLER_207_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8182_ _8182_/A _8995_/X vssd1 vssd1 vccd1 vccd1 _9528_/D sky130_fd_sc_hd__or2_1
X_7202_ _7487_/A _7491_/B vssd1 vssd1 vccd1 vccd1 _7202_/X sky130_fd_sc_hd__or2_2
X_5394_ _5389_/B _5379_/X _5392_/Y _5393_/Y _5364_/A vssd1 vssd1 vccd1 vccd1 _5395_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_132_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7133_ _9431_/X vssd1 vssd1 vccd1 vccd1 _7178_/B sky130_fd_sc_hd__buf_1
XFILLER_207_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7064_ _7064_/A vssd1 vssd1 vccd1 vccd1 _7073_/A sky130_fd_sc_hd__inv_2
X_6015_ _9853_/Q vssd1 vssd1 vccd1 vccd1 _7955_/A sky130_fd_sc_hd__inv_2
XFILLER_74_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7966_ _9634_/Q vssd1 vssd1 vccd1 vccd1 _7967_/A sky130_fd_sc_hd__inv_2
X_9705_ _9708_/CLK _9705_/D vssd1 vssd1 vccd1 vccd1 _9705_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7897_ _7897_/A _7897_/B vssd1 vssd1 vccd1 vccd1 _7902_/B sky130_fd_sc_hd__or2_2
X_6917_ _6742_/A _6742_/B _6743_/B vssd1 vssd1 vccd1 vccd1 _6917_/X sky130_fd_sc_hd__a21bo_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9636_ _9650_/CLK _9636_/D vssd1 vssd1 vccd1 vccd1 _9636_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_50_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6848_ _6845_/X _6847_/X _6845_/X _6847_/X vssd1 vssd1 vccd1 vccd1 _6848_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_210_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9567_ _9888_/CLK _9567_/D vssd1 vssd1 vccd1 vccd1 _9567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8518_ _9632_/Q _8580_/B _8545_/C _8517_/X vssd1 vssd1 vccd1 vccd1 _8518_/X sky130_fd_sc_hd__a31o_1
XPHY_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6779_ _6779_/A vssd1 vssd1 vccd1 vccd1 _6781_/A sky130_fd_sc_hd__inv_2
XFILLER_182_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9498_ _9497_/X _6981_/A _9507_/S vssd1 vssd1 vccd1 vccd1 _9498_/X sky130_fd_sc_hd__mux2_1
X_8449_ _8534_/A _9379_/X _8472_/A _8469_/B vssd1 vssd1 vccd1 vccd1 _8450_/B sky130_fd_sc_hd__o22a_1
XFILLER_184_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7820_ _9907_/Q _7815_/Y _7818_/X _7823_/B vssd1 vssd1 vccd1 vccd1 _7820_/X sky130_fd_sc_hd__o211a_1
XFILLER_76_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7751_ _7882_/A _9773_/Q _8123_/A _6371_/A _7750_/X vssd1 vssd1 vccd1 vccd1 _7752_/D
+ sky130_fd_sc_hd__o221a_1
X_4963_ input7/X input8/X _9038_/S vssd1 vssd1 vccd1 vccd1 _8047_/B sky130_fd_sc_hd__or3_4
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7682_ _7682_/A _7889_/A vssd1 vssd1 vccd1 vccd1 _7683_/B sky130_fd_sc_hd__or2_1
X_6702_ _9094_/X vssd1 vssd1 vccd1 vccd1 _6705_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9421_ _8888_/X _8886_/A _9490_/S vssd1 vssd1 vccd1 vccd1 _9421_/X sky130_fd_sc_hd__mux2_2
X_4894_ _5339_/A vssd1 vssd1 vccd1 vccd1 _5348_/B sky130_fd_sc_hd__inv_2
X_6633_ _6642_/A vssd1 vssd1 vccd1 vccd1 _6678_/A sky130_fd_sc_hd__buf_1
XFILLER_164_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater90 _9148_/S vssd1 vssd1 vccd1 vccd1 _9155_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_118_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9352_ _7055_/X _7632_/Y _9683_/Q vssd1 vssd1 vccd1 vccd1 _9352_/X sky130_fd_sc_hd__mux2_2
X_6564_ _6564_/A vssd1 vssd1 vccd1 vccd1 _6564_/X sky130_fd_sc_hd__clkbuf_2
X_6495_ _6304_/Y _6482_/X _6487_/X _6493_/X _6494_/Y vssd1 vssd1 vccd1 vccd1 _6495_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_145_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5515_ _9684_/Q vssd1 vssd1 vccd1 vccd1 _5515_/X sky130_fd_sc_hd__buf_2
X_8303_ _9544_/Q vssd1 vssd1 vccd1 vccd1 _8303_/Y sky130_fd_sc_hd__inv_2
X_9283_ _7843_/Y _9764_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9283_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8234_ _6335_/A _8232_/B _8232_/X vssd1 vssd1 vccd1 vccd1 _8234_/Y sky130_fd_sc_hd__a21boi_1
X_5446_ _6796_/C vssd1 vssd1 vccd1 vccd1 _6872_/A sky130_fd_sc_hd__clkbuf_2
X_8165_ _4788_/X _8099_/Y _9920_/Q _8100_/Y _8164_/X vssd1 vssd1 vccd1 vccd1 _8165_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_160_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5377_ _5372_/B _5356_/X _5376_/Y _5330_/A _5364_/X vssd1 vssd1 vccd1 vccd1 _5378_/A
+ sky130_fd_sc_hd__o32a_1
X_8096_ _9556_/Q _8084_/B _8085_/B vssd1 vssd1 vccd1 vccd1 _8096_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_141_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7116_ _7178_/A vssd1 vssd1 vccd1 vccd1 _7497_/A sky130_fd_sc_hd__buf_2
XFILLER_101_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7047_ _6945_/X _6952_/X _6945_/X _6952_/X vssd1 vssd1 vccd1 vccd1 _7064_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8998_ _8997_/X _9522_/Q _9155_/S vssd1 vssd1 vccd1 vccd1 _8998_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7949_ _7949_/A _9013_/S vssd1 vssd1 vccd1 vccd1 _7949_/Y sky130_fd_sc_hd__nor2_1
XPHY_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9619_ _9715_/CLK _9619_/D vssd1 vssd1 vccd1 vccd1 _9619_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5300_ _5295_/B _5224_/A _5299_/Y _5275_/A _5241_/A vssd1 vssd1 vccd1 vccd1 _5301_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6280_ _9590_/Q _6170_/A _8038_/A _6140_/A vssd1 vssd1 vccd1 vccd1 _6285_/A sky130_fd_sc_hd__a22o_1
XFILLER_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5231_ _9739_/Q vssd1 vssd1 vccd1 vccd1 _5244_/A sky130_fd_sc_hd__inv_2
X_5162_ _9775_/Q vssd1 vssd1 vccd1 vccd1 _5162_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_142_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5093_ _5214_/A vssd1 vssd1 vccd1 vccd1 _8177_/A sky130_fd_sc_hd__buf_2
XFILLER_84_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8921_ _8920_/A _8920_/B _8920_/Y vssd1 vssd1 vccd1 vccd1 _8921_/X sky130_fd_sc_hd__a21o_1
XFILLER_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8852_ _8774_/A _8851_/A _8775_/B _8851_/Y vssd1 vssd1 vccd1 vccd1 _8852_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8783_ _8810_/A _8810_/B _8810_/A _8810_/B vssd1 vssd1 vccd1 vccd1 _8783_/X sky130_fd_sc_hd__a2bb2o_1
X_7803_ _7803_/A _7803_/B vssd1 vssd1 vccd1 vccd1 _7807_/B sky130_fd_sc_hd__or2_4
XFILLER_64_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7734_ _7682_/A _6344_/Y _4812_/X _6429_/Y _7733_/X vssd1 vssd1 vccd1 vccd1 _7752_/A
+ sky130_fd_sc_hd__o221a_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5995_ _7941_/A _9638_/Q vssd1 vssd1 vccd1 vccd1 _5998_/A sky130_fd_sc_hd__nor2_1
X_4946_ _9120_/X _4943_/X _9857_/Q _4944_/X _4939_/X vssd1 vssd1 vccd1 vccd1 _9857_/D
+ sky130_fd_sc_hd__o221a_1
X_7665_ _7665_/A _7665_/B vssd1 vssd1 vccd1 vccd1 _7821_/A sky130_fd_sc_hd__or2_1
X_4877_ _9742_/Q _4870_/X _9890_/Q _4871_/X _4873_/X vssd1 vssd1 vccd1 vccd1 _9890_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9404_ _7999_/X _6094_/B _9504_/S vssd1 vssd1 vccd1 vccd1 _9404_/X sky130_fd_sc_hd__mux2_1
X_6616_ _6877_/A vssd1 vssd1 vccd1 vccd1 _6707_/A sky130_fd_sc_hd__buf_1
X_7596_ _7596_/A _7596_/B vssd1 vssd1 vccd1 vccd1 _7597_/B sky130_fd_sc_hd__or2_1
X_6547_ _6547_/A _6547_/B vssd1 vssd1 vccd1 vccd1 _6547_/Y sky130_fd_sc_hd__nor2_1
X_9335_ _5975_/X _5971_/A _9523_/Q vssd1 vssd1 vccd1 vccd1 _9335_/X sky130_fd_sc_hd__mux2_4
XFILLER_192_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6478_ _6478_/A vssd1 vssd1 vccd1 vccd1 _6478_/Y sky130_fd_sc_hd__inv_2
X_9266_ _9265_/X input17/X _9294_/S vssd1 vssd1 vccd1 vccd1 _9266_/X sky130_fd_sc_hd__mux2_1
X_9197_ _6540_/Y _9802_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9551_/D sky130_fd_sc_hd__mux2_1
X_8217_ _8213_/A _8219_/B _6349_/Y _8216_/Y vssd1 vssd1 vccd1 vccd1 _8217_/X sky130_fd_sc_hd__o22a_1
XFILLER_106_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5429_ _9343_/X vssd1 vssd1 vccd1 vccd1 _5431_/A sky130_fd_sc_hd__inv_2
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8148_ _7761_/X _8115_/X _8147_/Y vssd1 vssd1 vccd1 vccd1 _8148_/X sky130_fd_sc_hd__o21ba_1
XFILLER_87_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_1 _8955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8079_ _9551_/Q _8079_/B vssd1 vssd1 vccd1 vccd1 _8080_/B sky130_fd_sc_hd__or2_2
XFILLER_87_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4800_ _9298_/X _4796_/X _4798_/X _4799_/X _4791_/X vssd1 vssd1 vccd1 vccd1 _9918_/D
+ sky130_fd_sc_hd__o221a_1
X_5780_ _9661_/Q _5774_/X _5769_/X _7109_/A _5772_/X vssd1 vssd1 vccd1 vccd1 _9661_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_9_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7450_ _7374_/A _7374_/B _7376_/A vssd1 vssd1 vccd1 vccd1 _7450_/X sky130_fd_sc_hd__a21bo_1
X_6401_ _6549_/B vssd1 vssd1 vccd1 vccd1 _6401_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9120_ _9604_/Q input47/X _9667_/Q vssd1 vssd1 vccd1 vccd1 _9120_/X sky130_fd_sc_hd__mux2_1
X_7381_ _7407_/A _7400_/B _7400_/A _7398_/B vssd1 vssd1 vccd1 vccd1 _7381_/X sky130_fd_sc_hd__or4_4
XFILLER_127_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6332_ _9793_/Q vssd1 vssd1 vccd1 vccd1 _6456_/A sky130_fd_sc_hd__inv_2
X_6263_ _9587_/Q vssd1 vssd1 vccd1 vccd1 _8031_/A sky130_fd_sc_hd__inv_2
XFILLER_115_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9051_ _8010_/Y _9610_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9051_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5214_ _5214_/A vssd1 vssd1 vccd1 vccd1 _5214_/X sky130_fd_sc_hd__buf_2
X_8002_ _9418_/X _8002_/B vssd1 vssd1 vccd1 vccd1 _8002_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6194_ _7988_/A _6193_/X _6200_/A _6189_/X vssd1 vssd1 vccd1 vccd1 _6194_/Y sky130_fd_sc_hd__o22ai_1
X_5145_ _5045_/X _9780_/Q _5138_/A _9207_/X _5140_/X vssd1 vssd1 vccd1 vccd1 _9780_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5076_ _9805_/Q vssd1 vssd1 vccd1 vccd1 _6317_/C sky130_fd_sc_hd__inv_2
XFILLER_84_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8904_ _8904_/A _8904_/B vssd1 vssd1 vccd1 vccd1 _8904_/X sky130_fd_sc_hd__or2_1
XFILLER_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9884_ _9888_/CLK _9884_/D vssd1 vssd1 vccd1 vccd1 _9884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8835_ _8820_/X _8834_/X _8820_/X _8834_/X vssd1 vssd1 vccd1 vccd1 _8835_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8766_ _8955_/A _8766_/B _8766_/C vssd1 vssd1 vccd1 vccd1 _8766_/X sky130_fd_sc_hd__or3_2
X_5978_ _9849_/Q vssd1 vssd1 vccd1 vccd1 _7928_/A sky130_fd_sc_hd__inv_2
XFILLER_178_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8697_ _8385_/X _8406_/X _8385_/X _8406_/X vssd1 vssd1 vccd1 vccd1 _8698_/A sky130_fd_sc_hd__a2bb2o_1
X_7717_ _7713_/X _6331_/A _4798_/X _6349_/Y _7716_/X vssd1 vssd1 vccd1 vccd1 _7731_/B
+ sky130_fd_sc_hd__o221a_1
X_4929_ input5/X input4/X _4929_/C _4856_/C vssd1 vssd1 vccd1 vccd1 _5862_/A sky130_fd_sc_hd__or4b_4
XFILLER_178_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7648_ _7648_/A _7648_/B vssd1 vssd1 vccd1 vccd1 _7648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7579_ _7535_/X _7551_/X _7535_/X _7551_/X vssd1 vssd1 vccd1 vccd1 _7580_/A sky130_fd_sc_hd__a2bb2o_1
X_9318_ _9317_/X input35/X _9334_/S vssd1 vssd1 vccd1 vccd1 _9318_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9249_ _9248_/X _7804_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9249_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6950_ _6851_/A _6851_/B _6851_/X vssd1 vssd1 vccd1 vccd1 _6951_/B sky130_fd_sc_hd__a21bo_1
XFILLER_93_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5901_ _5903_/A _9139_/X vssd1 vssd1 vccd1 vccd1 _9608_/D sky130_fd_sc_hd__and2_1
XFILLER_81_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6881_ _6890_/B _6881_/B vssd1 vssd1 vccd1 vccd1 _6882_/A sky130_fd_sc_hd__or2_2
X_8620_ _8620_/A vssd1 vssd1 vccd1 vccd1 _8620_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5832_ _5832_/A vssd1 vssd1 vccd1 vccd1 _5832_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8551_ _8542_/X _8550_/Y _8542_/X _8550_/Y vssd1 vssd1 vccd1 vccd1 _8551_/X sky130_fd_sc_hd__a2bb2o_1
X_5763_ _5714_/X _5756_/X _5714_/X _5756_/X vssd1 vssd1 vccd1 vccd1 _7492_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7502_ _7502_/A _7502_/B vssd1 vssd1 vccd1 vccd1 _7503_/B sky130_fd_sc_hd__nor2_1
X_8482_ _8495_/A _8481_/B _8481_/X vssd1 vssd1 vccd1 vccd1 _8483_/B sky130_fd_sc_hd__a21bo_1
XFILLER_175_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5694_ _9672_/Q _5689_/X _9099_/X _5692_/X _5690_/X vssd1 vssd1 vccd1 vccd1 _9672_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_107_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7433_ _7306_/X _7376_/X _7306_/X _7376_/X vssd1 vssd1 vccd1 vccd1 _7433_/X sky130_fd_sc_hd__a2bb2o_1
X_7364_ _7362_/X _7363_/X _7362_/X _7363_/X vssd1 vssd1 vccd1 vccd1 _7364_/X sky130_fd_sc_hd__a2bb2o_1
X_6315_ _6315_/A _6315_/B _6315_/C _6315_/D vssd1 vssd1 vccd1 vccd1 _6315_/Y sky130_fd_sc_hd__nor4_2
X_9103_ _6050_/Y _6051_/Y _9896_/Q vssd1 vssd1 vccd1 vccd1 _9103_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9034_ _7982_/Y _9033_/X _9052_/S vssd1 vssd1 vccd1 vccd1 _9034_/X sky130_fd_sc_hd__mux2_1
X_7295_ _7278_/X _7279_/X _7278_/X _7279_/X vssd1 vssd1 vccd1 vccd1 _7296_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6246_ _8017_/A _6245_/X _8019_/A _6245_/X _6234_/B vssd1 vssd1 vccd1 vccd1 _6247_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_103_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6177_ _7965_/A _6197_/A _7973_/A _6135_/A vssd1 vssd1 vccd1 vccd1 _6177_/X sky130_fd_sc_hd__o22a_1
XFILLER_57_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5128_ _5128_/A vssd1 vssd1 vccd1 vccd1 _5128_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5059_ _5045_/X _6316_/C _5058_/Y _5050_/X vssd1 vssd1 vccd1 vccd1 _5060_/B sky130_fd_sc_hd__o22a_1
XFILLER_84_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9867_ _9874_/CLK _9867_/D vssd1 vssd1 vccd1 vccd1 _9867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8818_ _8959_/A _8955_/B vssd1 vssd1 vccd1 vccd1 _8818_/X sky130_fd_sc_hd__or2_1
XFILLER_111_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9798_ _9916_/CLK _9798_/D vssd1 vssd1 vccd1 vccd1 _9798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8749_ _8732_/X _8738_/X _8739_/X _8740_/X vssd1 vssd1 vccd1 vccd1 _8749_/X sky130_fd_sc_hd__o22a_1
XFILLER_40_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6100_ _9862_/Q vssd1 vssd1 vccd1 vccd1 _8003_/A sky130_fd_sc_hd__inv_2
XFILLER_140_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7080_ _7080_/A _7080_/B vssd1 vssd1 vccd1 vccd1 _7081_/B sky130_fd_sc_hd__or2_1
XFILLER_112_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6031_ _6031_/A vssd1 vssd1 vccd1 vccd1 _6031_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7982_ _8984_/X _7987_/B vssd1 vssd1 vccd1 vccd1 _7982_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9721_ _9893_/CLK _9721_/D vssd1 vssd1 vccd1 vccd1 _9721_/Q sky130_fd_sc_hd__dfxtp_1
X_6933_ _6929_/X _6930_/X _6929_/X _6930_/X vssd1 vssd1 vccd1 vccd1 _6933_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9652_ _9673_/CLK _9652_/D vssd1 vssd1 vccd1 vccd1 _9652_/Q sky130_fd_sc_hd__dfxtp_1
X_6864_ _6890_/B _6883_/B _6883_/A _6881_/B vssd1 vssd1 vccd1 vccd1 _6864_/X sky130_fd_sc_hd__or4_4
XFILLER_179_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8603_ _8603_/A _8603_/B vssd1 vssd1 vccd1 vccd1 _8650_/A sky130_fd_sc_hd__or2_1
X_5815_ _5815_/A _5815_/B _5862_/A _5815_/D vssd1 vssd1 vccd1 vccd1 _7911_/A sky130_fd_sc_hd__or4_4
XFILLER_22_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9583_ _9833_/CLK _9583_/D vssd1 vssd1 vccd1 vccd1 _9583_/Q sky130_fd_sc_hd__dfxtp_1
X_6795_ _6795_/A _6794_/X vssd1 vssd1 vccd1 vccd1 _6795_/X sky130_fd_sc_hd__or2b_1
XFILLER_210_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8534_ _8534_/A _9381_/X vssd1 vssd1 vccd1 vccd1 _8610_/C sky130_fd_sc_hd__or2_2
XFILLER_179_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5746_ _6567_/A _9654_/Q _5740_/Y _5745_/X vssd1 vssd1 vccd1 vccd1 _5746_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8465_ _8392_/X _8400_/X _8392_/X _8400_/X vssd1 vssd1 vccd1 vccd1 _8466_/A sky130_fd_sc_hd__a2bb2o_1
X_5677_ _9683_/Q _5671_/X _9110_/X _5676_/X _5674_/X vssd1 vssd1 vccd1 vccd1 _9683_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_175_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7416_ _7416_/A vssd1 vssd1 vccd1 vccd1 _7442_/A sky130_fd_sc_hd__inv_2
XFILLER_163_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8396_ _9685_/Q _6571_/Y _9685_/Q _6571_/Y vssd1 vssd1 vccd1 vccd1 _8396_/X sky130_fd_sc_hd__a2bb2o_1
X_7347_ _7347_/A _7347_/B vssd1 vssd1 vccd1 vccd1 _7348_/B sky130_fd_sc_hd__or2_2
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7278_ _7268_/X _7269_/X _7276_/X _7277_/X vssd1 vssd1 vccd1 vccd1 _7278_/X sky130_fd_sc_hd__o22a_1
XFILLER_131_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6229_ _6232_/B _6228_/Y _6232_/B _6228_/Y vssd1 vssd1 vccd1 vccd1 _6229_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9017_ _7943_/Y _9598_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9017_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9919_ _9923_/CLK _9919_/D vssd1 vssd1 vccd1 vccd1 _9919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput61 _9054_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_107_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput50 _9930_/Q vssd1 vssd1 vccd1 vccd1 io_irq sky130_fd_sc_hd__clkbuf_2
Xoutput72 _9064_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_110_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput83 _9515_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5600_ _5600_/A _5600_/B vssd1 vssd1 vccd1 vccd1 _5600_/Y sky130_fd_sc_hd__nor2_1
X_6580_ _6578_/A _6578_/B _6579_/Y vssd1 vssd1 vccd1 vccd1 _6580_/X sky130_fd_sc_hd__a21o_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5531_ _5595_/A _5595_/B vssd1 vssd1 vccd1 vccd1 _5594_/A sky130_fd_sc_hd__nand2_1
XFILLER_157_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8250_ _8191_/A _8191_/B _8231_/B vssd1 vssd1 vccd1 vccd1 _8250_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5462_ _9348_/X _9346_/X _5412_/Y _5475_/A vssd1 vssd1 vccd1 vccd1 _5471_/A sky130_fd_sc_hd__o22a_1
X_7201_ _7201_/A vssd1 vssd1 vccd1 vccd1 _7487_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_160_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8181_ _8182_/A _9444_/X vssd1 vssd1 vccd1 vccd1 _9527_/D sky130_fd_sc_hd__or2_1
X_5393_ _9719_/Q vssd1 vssd1 vccd1 vccd1 _5393_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7132_ _7223_/A vssd1 vssd1 vccd1 vccd1 _7494_/A sky130_fd_sc_hd__buf_2
XFILLER_140_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7063_ _7063_/A vssd1 vssd1 vccd1 vccd1 _7074_/A sky130_fd_sc_hd__inv_2
XFILLER_113_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6014_ _9853_/Q _6014_/B vssd1 vssd1 vccd1 vccd1 _6017_/A sky130_fd_sc_hd__nor2_1
XFILLER_100_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9704_ _9819_/CLK _9704_/D vssd1 vssd1 vccd1 vccd1 _9704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7965_ _7965_/A _9013_/S vssd1 vssd1 vccd1 vccd1 _7965_/Y sky130_fd_sc_hd__nor2_1
X_7896_ _7897_/A _7889_/Y _7683_/B vssd1 vssd1 vccd1 vccd1 _7896_/Y sky130_fd_sc_hd__o21ai_1
XPHY_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6916_ _6884_/X _6905_/X _6884_/X _6905_/X vssd1 vssd1 vccd1 vccd1 _6916_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9635_ _9828_/CLK _9635_/D vssd1 vssd1 vccd1 vccd1 _9635_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6847_ _6847_/A _6847_/B vssd1 vssd1 vccd1 vccd1 _6847_/X sky130_fd_sc_hd__or2_1
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6778_ _6761_/X _6762_/X _6761_/X _6762_/X vssd1 vssd1 vccd1 vccd1 _6779_/A sky130_fd_sc_hd__a2bb2o_1
X_9566_ _9888_/CLK _9566_/D vssd1 vssd1 vccd1 vccd1 _9566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8517_ _8875_/A _8626_/B _8776_/A _8543_/B vssd1 vssd1 vccd1 vccd1 _8517_/X sky130_fd_sc_hd__o22a_1
X_5729_ _9659_/Q vssd1 vssd1 vccd1 vccd1 _5729_/Y sky130_fd_sc_hd__inv_2
XFILLER_210_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9497_ _9496_/X _7491_/A _9506_/S vssd1 vssd1 vccd1 vccd1 _9497_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8448_ _9630_/Q _8580_/B _8472_/C vssd1 vssd1 vccd1 vccd1 _8499_/A sky130_fd_sc_hd__and3_1
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8379_ _9698_/Q _6598_/X _9698_/Q _6598_/X vssd1 vssd1 vccd1 vccd1 _8379_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_2_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7750_ _4835_/X _7748_/Y _8322_/A _5218_/X vssd1 vssd1 vccd1 vccd1 _7750_/X sky130_fd_sc_hd__o22a_1
XFILLER_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4962_ _4962_/A vssd1 vssd1 vccd1 vccd1 _9038_/S sky130_fd_sc_hd__clkbuf_4
X_7681_ _9924_/Q _7681_/B vssd1 vssd1 vccd1 vccd1 _7889_/A sky130_fd_sc_hd__or2_1
X_4893_ _9930_/Q _5048_/A vssd1 vssd1 vccd1 vccd1 _5339_/A sky130_fd_sc_hd__or2_2
X_6701_ _6701_/A _6700_/X vssd1 vssd1 vccd1 vccd1 _6701_/X sky130_fd_sc_hd__or2b_1
XFILLER_32_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9420_ _8932_/X _8930_/A _9490_/S vssd1 vssd1 vccd1 vccd1 _9420_/X sky130_fd_sc_hd__mux2_2
X_6632_ _6660_/A _6971_/B _6766_/A _6660_/B vssd1 vssd1 vccd1 vccd1 _6632_/X sky130_fd_sc_hd__or4_4
XFILLER_177_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater91 _9053_/S vssd1 vssd1 vccd1 vccd1 _9069_/S sky130_fd_sc_hd__buf_8
X_6563_ _6556_/A _6556_/B _6557_/B vssd1 vssd1 vccd1 vccd1 _6563_/X sky130_fd_sc_hd__a21bo_1
X_9351_ _7061_/A _7616_/X _9683_/Q vssd1 vssd1 vccd1 vccd1 _9351_/X sky130_fd_sc_hd__mux2_1
X_8302_ _8298_/Y _8302_/B _8302_/C vssd1 vssd1 vccd1 vccd1 _8377_/A sky130_fd_sc_hd__nand3b_1
X_5514_ _9627_/Q vssd1 vssd1 vccd1 vccd1 _8452_/A sky130_fd_sc_hd__inv_2
X_6494_ _6494_/A vssd1 vssd1 vccd1 vccd1 _6494_/Y sky130_fd_sc_hd__inv_2
X_9282_ _9281_/X input22/X _9282_/S vssd1 vssd1 vccd1 vccd1 _9282_/X sky130_fd_sc_hd__mux2_1
X_8233_ _9761_/Q _8232_/X _8229_/X vssd1 vssd1 vccd1 vccd1 _8233_/Y sky130_fd_sc_hd__a21boi_1
X_5445_ _7334_/B vssd1 vssd1 vccd1 vccd1 _7389_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_172_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8164_ _4794_/A _8101_/Y _9920_/Q _8100_/Y _8163_/X vssd1 vssd1 vccd1 vccd1 _8164_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_160_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5376_ _9723_/Q _5376_/B vssd1 vssd1 vccd1 vccd1 _5376_/Y sky130_fd_sc_hd__nor2_1
X_7115_ _7290_/A vssd1 vssd1 vccd1 vccd1 _7178_/A sky130_fd_sc_hd__buf_1
X_8095_ _9557_/Q _8085_/B _8093_/Y vssd1 vssd1 vccd1 vccd1 _8095_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_99_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7046_ _6954_/A _6954_/B _6954_/Y vssd1 vssd1 vccd1 vccd1 _7063_/A sky130_fd_sc_hd__o21ai_1
XFILLER_170_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8997_ _9522_/Q _5039_/A _8999_/S vssd1 vssd1 vccd1 vccd1 _8997_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7948_ _9489_/X _7956_/B vssd1 vssd1 vccd1 vccd1 _7948_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7879_ _7879_/A vssd1 vssd1 vccd1 vccd1 _7879_/Y sky130_fd_sc_hd__inv_2
XPHY_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9618_ _9656_/CLK _9618_/D vssd1 vssd1 vccd1 vccd1 _9618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9549_ _9923_/CLK _9549_/D vssd1 vssd1 vccd1 vccd1 _9549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5230_ _9740_/Q vssd1 vssd1 vccd1 vccd1 _5245_/A sky130_fd_sc_hd__inv_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5161_ _8200_/A _5155_/X input36/X _5157_/X _5153_/X vssd1 vssd1 vccd1 vccd1 _9776_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5092_ _5092_/A _5092_/B vssd1 vssd1 vccd1 vccd1 _9802_/D sky130_fd_sc_hd__nor2_1
X_8920_ _8920_/A _8920_/B vssd1 vssd1 vccd1 vccd1 _8920_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8851_ _8851_/A vssd1 vssd1 vccd1 vccd1 _8851_/Y sky130_fd_sc_hd__inv_2
X_8782_ _8781_/A _8781_/B _8811_/A vssd1 vssd1 vccd1 vccd1 _8810_/B sky130_fd_sc_hd__a21oi_1
X_7802_ _7803_/A _7795_/Y _7661_/B vssd1 vssd1 vccd1 vccd1 _7802_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5994_ _9851_/Q vssd1 vssd1 vccd1 vccd1 _7941_/A sky130_fd_sc_hd__inv_2
XFILLER_169_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7733_ _7696_/X _5198_/X _7788_/A _8183_/B vssd1 vssd1 vccd1 vccd1 _7733_/X sky130_fd_sc_hd__o2bb2a_1
X_4945_ _9121_/X _4943_/X _9858_/Q _4944_/X _4939_/X vssd1 vssd1 vccd1 vccd1 _9858_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7664_ _9907_/Q _7812_/A vssd1 vssd1 vccd1 vccd1 _7665_/B sky130_fd_sc_hd__or2_2
X_4876_ _9743_/Q _4870_/X _9891_/Q _4871_/X _4873_/X vssd1 vssd1 vccd1 vccd1 _9891_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9403_ _8556_/X _8554_/A _9490_/S vssd1 vssd1 vccd1 vccd1 _9403_/X sky130_fd_sc_hd__mux2_2
X_6615_ _9616_/Q vssd1 vssd1 vccd1 vccd1 _6877_/A sky130_fd_sc_hd__inv_2
X_7595_ _7595_/A _7595_/B vssd1 vssd1 vccd1 vccd1 _7596_/B sky130_fd_sc_hd__or2_1
X_9334_ _9333_/X input40/X _9334_/S vssd1 vssd1 vccd1 vccd1 _9334_/X sky130_fd_sc_hd__mux2_1
X_6546_ _6547_/A _6546_/B vssd1 vssd1 vccd1 vccd1 _6546_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6477_ _6309_/Y _6475_/X _9785_/Q _6519_/B vssd1 vssd1 vccd1 vccd1 _6478_/A sky130_fd_sc_hd__a2bb2o_1
X_9265_ _9264_/X _7820_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9265_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9196_ _6539_/Y _9801_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9550_/D sky130_fd_sc_hd__mux2_1
X_8216_ _9768_/Q _8216_/B vssd1 vssd1 vccd1 vccd1 _8216_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5428_ _9337_/X _9336_/X _9337_/X _9336_/X vssd1 vssd1 vccd1 vccd1 _5428_/X sky130_fd_sc_hd__a2bb2o_2
X_8147_ _7696_/X _8116_/X _8146_/X vssd1 vssd1 vccd1 vccd1 _8147_/Y sky130_fd_sc_hd__a21oi_1
X_5359_ _5353_/B _5356_/X _5358_/Y _5334_/A _5349_/X vssd1 vssd1 vccd1 vccd1 _5360_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8078_ _9550_/Q _8103_/A vssd1 vssd1 vccd1 vccd1 _8079_/B sky130_fd_sc_hd__or2_2
XINSDIODE2_2 _8047_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7029_ _6941_/X _6954_/Y _6955_/X _6957_/A vssd1 vssd1 vccd1 vccd1 _7030_/B sky130_fd_sc_hd__a31o_1
XFILLER_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6400_ _9778_/Q _8197_/A _6397_/Y vssd1 vssd1 vccd1 vccd1 _6549_/B sky130_fd_sc_hd__a21oi_2
XFILLER_147_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7380_ _7407_/A _7400_/B _7384_/C _7398_/B vssd1 vssd1 vccd1 vccd1 _7382_/A sky130_fd_sc_hd__o22a_1
XFILLER_134_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6331_ _6331_/A vssd1 vssd1 vccd1 vccd1 _6331_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6262_ _6265_/D _6261_/Y _6265_/D _6261_/Y vssd1 vssd1 vccd1 vccd1 _6262_/X sky130_fd_sc_hd__a2bb2o_1
X_9050_ _8007_/Y _9049_/X _9053_/S vssd1 vssd1 vccd1 vccd1 _9050_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6193_ _6193_/A vssd1 vssd1 vccd1 vccd1 _6193_/X sky130_fd_sc_hd__buf_4
X_5213_ _9751_/Q vssd1 vssd1 vccd1 vccd1 _8183_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8001_ _8001_/A _8010_/B vssd1 vssd1 vccd1 vccd1 _8001_/Y sky130_fd_sc_hd__nor2_1
X_5144_ _5045_/X _9781_/Q _5138_/X _9208_/X _5140_/X vssd1 vssd1 vccd1 vccd1 _9781_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5075_ _5092_/A _5075_/B vssd1 vssd1 vccd1 vccd1 _9806_/D sky130_fd_sc_hd__nor2_1
XFILLER_96_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8903_ _8903_/A vssd1 vssd1 vccd1 vccd1 _8903_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9883_ _9895_/CLK _9883_/D vssd1 vssd1 vccd1 vccd1 _9883_/Q sky130_fd_sc_hd__dfxtp_1
X_8834_ _8903_/A _8833_/B _8833_/Y vssd1 vssd1 vccd1 vccd1 _8834_/X sky130_fd_sc_hd__a21o_1
XFILLER_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8765_ _8765_/A vssd1 vssd1 vccd1 vccd1 _8765_/Y sky130_fd_sc_hd__inv_2
X_5977_ _7971_/A vssd1 vssd1 vccd1 vccd1 _9013_/S sky130_fd_sc_hd__buf_2
XFILLER_25_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8696_ _8695_/A _8695_/B _8743_/A vssd1 vssd1 vccd1 vccd1 _8696_/X sky130_fd_sc_hd__a21bo_1
X_7716_ _7715_/X _9763_/Q _4814_/X _6331_/Y vssd1 vssd1 vccd1 vccd1 _7716_/X sky130_fd_sc_hd__o22a_1
XFILLER_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4928_ input3/X input6/X vssd1 vssd1 vccd1 vccd1 _4931_/C sky130_fd_sc_hd__nand2_1
XFILLER_178_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7647_ _7647_/A _7648_/B vssd1 vssd1 vccd1 vccd1 _7647_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _4859_/A vssd1 vssd1 vccd1 vccd1 _8999_/S sky130_fd_sc_hd__inv_2
XFILLER_165_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7578_ _7578_/A vssd1 vssd1 vccd1 vccd1 _7604_/A sky130_fd_sc_hd__inv_2
X_9317_ _9316_/X _7894_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9317_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6529_ _6529_/A _6529_/B vssd1 vssd1 vccd1 vccd1 _6529_/Y sky130_fd_sc_hd__nor2_1
X_9248_ _9754_/Q _9247_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9248_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9179_ _9178_/X _9784_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9533_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5900_ _5903_/A _9140_/X vssd1 vssd1 vccd1 vccd1 _9609_/D sky130_fd_sc_hd__and2_1
XFILLER_207_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6880_ _6865_/X _6867_/X _6878_/X _6879_/X vssd1 vssd1 vccd1 vccd1 _6880_/X sky130_fd_sc_hd__o22a_1
XFILLER_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5831_ _9643_/Q _5824_/X input46/X _5825_/X _5830_/X vssd1 vssd1 vccd1 vccd1 _9643_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_201_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8550_ _8626_/C _8549_/B _8591_/A vssd1 vssd1 vccd1 vccd1 _8550_/Y sky130_fd_sc_hd__o21ai_2
X_5762_ _9666_/Q _5697_/X _5570_/X _7492_/D _5698_/X vssd1 vssd1 vccd1 vccd1 _9666_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7501_ _7186_/A _7192_/A _7186_/Y vssd1 vssd1 vccd1 vccd1 _7501_/X sky130_fd_sc_hd__a21o_1
X_8481_ _8495_/A _8481_/B vssd1 vssd1 vccd1 vccd1 _8481_/X sky130_fd_sc_hd__or2_1
XFILLER_175_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5693_ _6556_/A _5689_/X _9100_/X _5692_/X _5690_/X vssd1 vssd1 vccd1 vccd1 _9673_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7432_ _7401_/X _7422_/X _7401_/X _7422_/X vssd1 vssd1 vccd1 vccd1 _7432_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_162_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7363_ _7348_/B _7350_/B _7350_/X vssd1 vssd1 vccd1 vccd1 _7363_/X sky130_fd_sc_hd__o21a_1
XFILLER_162_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6314_ _9791_/Q _9790_/Q _9789_/Q _9788_/Q vssd1 vssd1 vccd1 vccd1 _6315_/D sky130_fd_sc_hd__or4_4
XFILLER_115_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9102_ _6038_/X _6040_/X _9896_/Q vssd1 vssd1 vccd1 vccd1 _9102_/X sky130_fd_sc_hd__mux2_1
X_7294_ _7289_/X _7293_/X _7289_/X _7293_/X vssd1 vssd1 vccd1 vccd1 _7294_/X sky130_fd_sc_hd__a2bb2o_1
X_6245_ _6245_/A vssd1 vssd1 vccd1 vccd1 _6245_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9033_ _7983_/Y _9604_/Q _9051_/S vssd1 vssd1 vccd1 vccd1 _9033_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6176_ _6176_/A _6159_/X vssd1 vssd1 vccd1 vccd1 _6176_/X sky130_fd_sc_hd__or2b_1
X_5127_ _4743_/X _9792_/Q _5121_/X _9219_/X _5124_/X vssd1 vssd1 vccd1 vccd1 _9792_/D
+ sky130_fd_sc_hd__o221a_1
X_5058_ _9841_/Q vssd1 vssd1 vccd1 vccd1 _5058_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9866_ _9874_/CLK _9866_/D vssd1 vssd1 vccd1 vccd1 _9866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8817_ _8875_/D vssd1 vssd1 vccd1 vccd1 _8955_/B sky130_fd_sc_hd__clkbuf_2
X_9797_ _9916_/CLK _9797_/D vssd1 vssd1 vccd1 vccd1 _9797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8748_ _8747_/A _8747_/B _8797_/A vssd1 vssd1 vccd1 vccd1 _8748_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_111_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8679_ _8667_/X _8678_/X _8667_/X _8678_/X vssd1 vssd1 vccd1 vccd1 _8679_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6030_ _7955_/A _9640_/Q _6017_/A _6021_/X vssd1 vssd1 vccd1 vccd1 _6031_/A sky130_fd_sc_hd__o22a_1
XFILLER_98_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7981_ _7981_/A _7981_/B vssd1 vssd1 vccd1 vccd1 _7981_/X sky130_fd_sc_hd__or2_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9720_ _9874_/CLK _9720_/D vssd1 vssd1 vccd1 vccd1 _9720_/Q sky130_fd_sc_hd__dfxtp_1
X_6932_ _6921_/X _6931_/X _6921_/X _6931_/X vssd1 vssd1 vccd1 vccd1 _6932_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_207_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9651_ _9715_/CLK _9651_/D vssd1 vssd1 vccd1 vccd1 _9651_/Q sky130_fd_sc_hd__dfxtp_1
X_6863_ _6890_/B _6883_/B _6867_/D _6881_/B vssd1 vssd1 vccd1 vccd1 _6865_/A sky130_fd_sc_hd__o22a_1
XFILLER_34_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8602_ _8602_/A vssd1 vssd1 vccd1 vccd1 _8603_/B sky130_fd_sc_hd__inv_2
X_5814_ _9651_/Q _5557_/X _4900_/X _7321_/D _5809_/X vssd1 vssd1 vccd1 vccd1 _9651_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_34_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9582_ _9833_/CLK _9582_/D vssd1 vssd1 vccd1 vccd1 _9582_/Q sky130_fd_sc_hd__dfxtp_1
X_6794_ _6821_/B _6868_/B _6796_/D _6862_/A vssd1 vssd1 vccd1 vccd1 _6794_/X sky130_fd_sc_hd__or4_4
XFILLER_210_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8533_ _8530_/X _8532_/X _8530_/X _8532_/X vssd1 vssd1 vccd1 vccd1 _8533_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_148_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5745_ _9670_/Q _9653_/Q _5741_/Y _5744_/Y vssd1 vssd1 vccd1 vccd1 _5745_/X sky130_fd_sc_hd__o2bb2a_1
X_8464_ _8463_/A _8463_/B _8486_/A vssd1 vssd1 vccd1 vccd1 _8464_/X sky130_fd_sc_hd__a21bo_1
XFILLER_175_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5676_ _5692_/A vssd1 vssd1 vccd1 vccd1 _5676_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7415_ _7415_/A _7421_/A vssd1 vssd1 vccd1 vccd1 _7415_/Y sky130_fd_sc_hd__nor2_1
XFILLER_190_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8395_ _9686_/Q _6569_/Y _9686_/Q _6569_/Y vssd1 vssd1 vccd1 vccd1 _8432_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_190_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7346_ _7346_/A _7346_/B vssd1 vssd1 vccd1 vccd1 _7347_/B sky130_fd_sc_hd__or2_1
X_7277_ _7487_/C _9469_/X _7277_/C vssd1 vssd1 vccd1 vccd1 _7277_/X sky130_fd_sc_hd__or3_1
X_9016_ _9015_/X _9751_/Q _9481_/S vssd1 vssd1 vccd1 vccd1 _9016_/X sky130_fd_sc_hd__mux2_2
X_6228_ _8013_/A _6143_/X _6232_/A vssd1 vssd1 vccd1 vccd1 _6228_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6159_ _7965_/A _6148_/X _9569_/Q _6165_/A vssd1 vssd1 vccd1 vccd1 _6159_/X sky130_fd_sc_hd__o22a_1
XFILLER_85_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9918_ _9923_/CLK _9918_/D vssd1 vssd1 vccd1 vccd1 _9918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9849_ _9879_/CLK _9849_/D vssd1 vssd1 vccd1 vccd1 _9849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput51 _9562_/Q vssd1 vssd1 vccd1 vccd1 io_pwm_h sky130_fd_sc_hd__clkbuf_2
XFILLER_122_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput73 _9065_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput62 _9055_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_110_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput84 _9032_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_163_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5530_ _9416_/X _5499_/X _5599_/A vssd1 vssd1 vccd1 vccd1 _5595_/B sky130_fd_sc_hd__o21ai_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5461_ _9360_/X _9356_/X _5415_/Y _5479_/A vssd1 vssd1 vccd1 vccd1 _5475_/A sky130_fd_sc_hd__o22a_1
XFILLER_172_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7200_ _7200_/A _7200_/B vssd1 vssd1 vccd1 vccd1 _7204_/A sky130_fd_sc_hd__or2_1
XFILLER_145_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8180_ _8182_/A _9445_/X vssd1 vssd1 vccd1 vccd1 _9526_/D sky130_fd_sc_hd__or2_1
X_5392_ _9719_/Q _5392_/B vssd1 vssd1 vccd1 vccd1 _5392_/Y sky130_fd_sc_hd__nor2_1
XFILLER_207_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7131_ _7385_/A vssd1 vssd1 vccd1 vccd1 _7223_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_207_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7062_ _7062_/A vssd1 vssd1 vccd1 vccd1 _7075_/A sky130_fd_sc_hd__inv_2
XFILLER_140_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6013_ _9640_/Q vssd1 vssd1 vccd1 vccd1 _6014_/B sky130_fd_sc_hd__inv_2
XFILLER_100_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7964_ _8978_/X _7987_/B vssd1 vssd1 vccd1 vccd1 _7964_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9703_ _9708_/CLK _9703_/D vssd1 vssd1 vccd1 vccd1 _9703_/Q sky130_fd_sc_hd__dfxtp_1
X_6915_ _6789_/X _6859_/X _6789_/X _6859_/X vssd1 vssd1 vccd1 vccd1 _6915_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7895_ _7895_/A vssd1 vssd1 vccd1 vccd1 _7897_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9634_ _9634_/CLK _9634_/D vssd1 vssd1 vccd1 vccd1 _9634_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6846_ _6846_/A _6846_/B vssd1 vssd1 vccd1 vccd1 _6847_/B sky130_fd_sc_hd__nor2_1
XFILLER_195_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6777_ _6772_/X _6776_/X _6772_/X _6776_/X vssd1 vssd1 vccd1 vccd1 _6777_/X sky130_fd_sc_hd__a2bb2o_2
X_9565_ _9888_/CLK _9565_/D vssd1 vssd1 vccd1 vccd1 _9565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8516_ _8516_/A vssd1 vssd1 vccd1 vccd1 _8545_/C sky130_fd_sc_hd__inv_2
XFILLER_148_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5728_ _9676_/Q vssd1 vssd1 vccd1 vccd1 _6582_/A sky130_fd_sc_hd__inv_2
XFILLER_136_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9496_ _9495_/X _8942_/A _9505_/S vssd1 vssd1 vccd1 vccd1 _9496_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8447_ _8445_/Y _8444_/X _8467_/A vssd1 vssd1 vccd1 vccd1 _8447_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_108_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5659_ _9673_/Q vssd1 vssd1 vccd1 vccd1 _6556_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_190_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8378_ _8378_/A _9052_/S _9038_/S vssd1 vssd1 vccd1 vccd1 _8378_/X sky130_fd_sc_hd__or3b_4
XFILLER_117_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7329_ _7334_/A _7379_/A vssd1 vssd1 vccd1 vccd1 _7330_/A sky130_fd_sc_hd__or2_2
XFILLER_117_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4961_ _5815_/D _5147_/A vssd1 vssd1 vccd1 vccd1 _4962_/A sky130_fd_sc_hd__or2_1
XFILLER_64_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7680_ _7680_/A _7879_/A vssd1 vssd1 vccd1 vccd1 _7681_/B sky130_fd_sc_hd__or2_1
X_4892_ _9929_/Q vssd1 vssd1 vccd1 vccd1 _5048_/A sky130_fd_sc_hd__inv_2
X_6700_ _6971_/A _6766_/B _7005_/A _6721_/B vssd1 vssd1 vccd1 vccd1 _6700_/X sky130_fd_sc_hd__or4_4
X_6631_ _6631_/A _6630_/X vssd1 vssd1 vccd1 vccd1 _6631_/X sky130_fd_sc_hd__or2b_1
XFILLER_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_9350_ _5467_/A _5467_/B _9350_/S vssd1 vssd1 vccd1 vccd1 _9350_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8301_ _8301_/A _8301_/B vssd1 vssd1 vccd1 vccd1 _8302_/C sky130_fd_sc_hd__nand2_1
XFILLER_145_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6562_ _6561_/A _6557_/B _6558_/B vssd1 vssd1 vccd1 vccd1 _6562_/X sky130_fd_sc_hd__a21bo_1
Xrepeater92 _9038_/S vssd1 vssd1 vccd1 vccd1 _9053_/S sky130_fd_sc_hd__buf_8
X_6493_ _9781_/Q _6329_/A _9780_/Q _6324_/A _6485_/X vssd1 vssd1 vccd1 vccd1 _6493_/X
+ sky130_fd_sc_hd__a221o_1
X_9281_ _9280_/X _7842_/Y _9526_/Q vssd1 vssd1 vccd1 vccd1 _9281_/X sky130_fd_sc_hd__mux2_1
X_5513_ _5513_/A _5450_/X vssd1 vssd1 vccd1 vccd1 _5627_/A sky130_fd_sc_hd__or2b_4
XFILLER_133_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8232_ _9760_/Q _8232_/B vssd1 vssd1 vccd1 vccd1 _8232_/X sky130_fd_sc_hd__or2_1
X_5444_ _7321_/D vssd1 vssd1 vccd1 vccd1 _7334_/B sky130_fd_sc_hd__inv_2
X_8163_ _4794_/A _8101_/Y _4798_/A _8104_/X _8162_/X vssd1 vssd1 vccd1 vccd1 _8163_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5375_ _5375_/A vssd1 vssd1 vccd1 vccd1 _5376_/B sky130_fd_sc_hd__inv_2
X_7114_ _7311_/A vssd1 vssd1 vccd1 vccd1 _7290_/A sky130_fd_sc_hd__buf_1
X_8094_ _8092_/Y _8093_/Y _8089_/B vssd1 vssd1 vccd1 vccd1 _8094_/X sky130_fd_sc_hd__o21a_1
XFILLER_101_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7045_ _7030_/A _7030_/B _7030_/X vssd1 vssd1 vccd1 vccd1 _7062_/A sky130_fd_sc_hd__a21bo_1
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8996_ _9525_/D _5041_/A _9445_/S vssd1 vssd1 vccd1 vccd1 _8996_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7947_ _7947_/A _9503_/S vssd1 vssd1 vccd1 vccd1 _7947_/X sky130_fd_sc_hd__or2_1
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7878_ _4788_/X _7874_/Y _7860_/X _7882_/B vssd1 vssd1 vccd1 vccd1 _7878_/X sky130_fd_sc_hd__o211a_1
XPHY_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_9617_ _9656_/CLK _9617_/D vssd1 vssd1 vccd1 vccd1 _9617_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6829_ _6829_/A _6835_/A vssd1 vssd1 vccd1 vccd1 _6829_/Y sky130_fd_sc_hd__nor2_1
XFILLER_195_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9548_ _9916_/CLK _9548_/D vssd1 vssd1 vccd1 vccd1 _9548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9479_ _9478_/X _6342_/Y _9481_/S vssd1 vssd1 vccd1 vccd1 _9479_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5160_ _9776_/Q vssd1 vssd1 vccd1 vccd1 _8200_/A sky130_fd_sc_hd__buf_2
XFILLER_96_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5091_ _5084_/X _6318_/B _5090_/Y _5073_/X vssd1 vssd1 vccd1 vccd1 _5092_/B sky130_fd_sc_hd__o22a_1
XFILLER_96_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8850_ _5843_/X _8656_/X _8893_/C _8849_/X vssd1 vssd1 vccd1 vccd1 _8851_/A sky130_fd_sc_hd__a31o_1
XFILLER_76_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8781_ _8781_/A _8781_/B vssd1 vssd1 vccd1 vccd1 _8811_/A sky130_fd_sc_hd__nor2_2
X_7801_ _7801_/A vssd1 vssd1 vccd1 vccd1 _7803_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_91_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5993_ _5989_/A _5992_/A _5987_/A _5992_/Y vssd1 vssd1 vccd1 vccd1 _5993_/X sky130_fd_sc_hd__o22a_1
XFILLER_64_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7732_ _9900_/Q vssd1 vssd1 vccd1 vccd1 _7788_/A sky130_fd_sc_hd__inv_2
X_4944_ _4952_/A vssd1 vssd1 vccd1 vccd1 _4944_/X sky130_fd_sc_hd__buf_1
XFILLER_24_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7663_ _9906_/Q _7663_/B vssd1 vssd1 vccd1 vccd1 _7812_/A sky130_fd_sc_hd__or2_1
X_9402_ _9401_/X _7005_/A _9507_/S vssd1 vssd1 vccd1 vccd1 _9402_/X sky130_fd_sc_hd__mux2_1
X_4875_ _9744_/Q _4870_/X _9892_/Q _4871_/X _4873_/X vssd1 vssd1 vccd1 vccd1 _9892_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_165_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6614_ _9617_/Q _6610_/Y _5890_/X _6612_/Y _6613_/X vssd1 vssd1 vccd1 vccd1 _6622_/A
+ sky130_fd_sc_hd__a41o_1
XFILLER_20_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7594_ _7594_/A _7594_/B vssd1 vssd1 vccd1 vccd1 _7595_/B sky130_fd_sc_hd__or2_1
X_9333_ _9332_/X _7910_/X _9526_/Q vssd1 vssd1 vccd1 vccd1 _9333_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6545_ _6547_/A _6545_/B vssd1 vssd1 vccd1 vccd1 _6545_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9264_ _9758_/Q _9263_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9264_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6476_ _6371_/A _6371_/B _6372_/B vssd1 vssd1 vccd1 vccd1 _6519_/B sky130_fd_sc_hd__o21a_1
XFILLER_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8215_ _8215_/A _8219_/B vssd1 vssd1 vccd1 vccd1 _8216_/B sky130_fd_sc_hd__or2_2
XFILLER_106_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_9195_ _6538_/Y _9800_/Q _9206_/S vssd1 vssd1 vccd1 vccd1 _9549_/D sky130_fd_sc_hd__mux2_1
X_5427_ _9364_/X _9362_/X _9364_/X _9362_/X vssd1 vssd1 vccd1 vccd1 _5427_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_160_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8146_ _7823_/A _8116_/X _8145_/X vssd1 vssd1 vccd1 vccd1 _8146_/X sky130_fd_sc_hd__o21a_1
X_5358_ _9727_/Q _5358_/B vssd1 vssd1 vccd1 vccd1 _5358_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8077_ _9549_/Q _8077_/B vssd1 vssd1 vccd1 vccd1 _8103_/A sky130_fd_sc_hd__or2_1
XINSDIODE2_3 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5289_ _5289_/A vssd1 vssd1 vccd1 vccd1 _9739_/D sky130_fd_sc_hd__inv_2
X_7028_ _7025_/X _7027_/X _7025_/X _7027_/X vssd1 vssd1 vccd1 vccd1 _7028_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8979_ _6340_/Y _7769_/Y _9480_/S vssd1 vssd1 vccd1 vccd1 _8979_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6330_ _9794_/Q vssd1 vssd1 vccd1 vccd1 _6330_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6261_ _8027_/A _6193_/X _6265_/C _6257_/X vssd1 vssd1 vccd1 vccd1 _6261_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_142_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5212_ _4978_/X _5203_/X _9752_/Q _5205_/X _5206_/X vssd1 vssd1 vccd1 vccd1 _9752_/D
+ sky130_fd_sc_hd__a221o_1
X_8000_ _9407_/X _8009_/B vssd1 vssd1 vccd1 vccd1 _8000_/Y sky130_fd_sc_hd__nor2_1
X_6192_ _9574_/Q _6167_/A _7993_/A _6137_/A vssd1 vssd1 vccd1 vccd1 _6200_/B sky130_fd_sc_hd__a22o_1
X_5143_ _5136_/X _9782_/Q _5138_/X _9209_/X _5140_/X vssd1 vssd1 vccd1 vccd1 _9782_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_111_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5074_ _5061_/X _6317_/B _5072_/Y _5073_/X vssd1 vssd1 vccd1 vccd1 _5075_/B sky130_fd_sc_hd__o22a_1
XFILLER_56_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8902_ _8900_/X _8901_/X _8900_/X _8901_/X vssd1 vssd1 vccd1 vccd1 _8902_/X sky130_fd_sc_hd__a2bb2o_1
X_9882_ _9895_/CLK _9882_/D vssd1 vssd1 vccd1 vccd1 _9882_/Q sky130_fd_sc_hd__dfxtp_1
X_8833_ _8903_/A _8833_/B vssd1 vssd1 vccd1 vccd1 _8833_/Y sky130_fd_sc_hd__nor2_1
XFILLER_197_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_8764_ _8728_/X _8729_/X _8730_/X _8731_/X vssd1 vssd1 vccd1 vccd1 _8765_/A sky130_fd_sc_hd__o22a_1
X_5976_ _5976_/A vssd1 vssd1 vccd1 vccd1 _7971_/A sky130_fd_sc_hd__inv_2
XFILLER_12_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8695_ _8695_/A _8695_/B vssd1 vssd1 vccd1 vccd1 _8743_/A sky130_fd_sc_hd__or2_1
X_7715_ _7840_/A vssd1 vssd1 vccd1 vccd1 _7715_/X sky130_fd_sc_hd__buf_2
XFILLER_33_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4927_ input7/X vssd1 vssd1 vccd1 vccd1 _5815_/A sky130_fd_sc_hd__inv_2
XFILLER_138_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7646_ _7646_/A _7648_/B vssd1 vssd1 vccd1 vccd1 _7646_/Y sky130_fd_sc_hd__nor2_1
X_4858_ _5816_/A _5976_/A vssd1 vssd1 vccd1 vccd1 _4859_/A sky130_fd_sc_hd__or2_1
XFILLER_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9316_ _9775_/Q _9315_/X _9525_/Q vssd1 vssd1 vccd1 vccd1 _9316_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4789_ _9306_/X _4782_/X _4788_/X _4784_/X _4778_/X vssd1 vssd1 vccd1 vccd1 _9921_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_109_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7577_ _7577_/A vssd1 vssd1 vccd1 vccd1 _7577_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_106_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6528_ _6529_/A _6528_/B vssd1 vssd1 vccd1 vccd1 _6528_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_9247_ _7802_/Y _9754_/Q _9291_/S vssd1 vssd1 vccd1 vccd1 _9247_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6459_ _9794_/Q _6531_/B vssd1 vssd1 vccd1 vccd1 _6463_/C sky130_fd_sc_hd__and2_1
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9178_ _9847_/Q _6475_/X _9178_/S vssd1 vssd1 vccd1 vccd1 _9178_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8129_ _8184_/A _9531_/Q _8053_/Y vssd1 vssd1 vccd1 vccd1 _8129_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5830_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5830_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5761_ _9475_/S vssd1 vssd1 vccd1 vccd1 _7492_/D sky130_fd_sc_hd__inv_2
X_8480_ _8479_/A _8479_/B _8479_/Y vssd1 vssd1 vccd1 vccd1 _8481_/B sky130_fd_sc_hd__a21o_1
XFILLER_15_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7500_ _7500_/A _7500_/B vssd1 vssd1 vccd1 vccd1 _7500_/X sky130_fd_sc_hd__or2_1
XFILLER_30_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5692_ _5692_/A vssd1 vssd1 vccd1 vccd1 _5692_/X sky130_fd_sc_hd__clkbuf_2
X_7431_ _7424_/X _7425_/X _7424_/X _7425_/X vssd1 vssd1 vccd1 vccd1 _7477_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7362_ _7352_/A _7352_/B _7352_/Y vssd1 vssd1 vccd1 vccd1 _7362_/X sky130_fd_sc_hd__a21o_1
XFILLER_143_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6313_ _9787_/Q _9786_/Q _9785_/Q vssd1 vssd1 vccd1 vccd1 _6315_/C sky130_fd_sc_hd__or3_1
X_9101_ _6029_/X _6032_/X _9896_/Q vssd1 vssd1 vccd1 vccd1 _9101_/X sky130_fd_sc_hd__mux2_1
X_7293_ _7283_/C _7292_/A _7282_/A _7292_/Y vssd1 vssd1 vccd1 vccd1 _7293_/X sky130_fd_sc_hd__a22o_1
X_6244_ _6244_/A _6244_/B _6244_/C vssd1 vssd1 vccd1 vccd1 _6247_/A sky130_fd_sc_hd__or3_4
X_9032_ _7980_/Y _9031_/X _9038_/S vssd1 vssd1 vccd1 vccd1 _9032_/X sky130_fd_sc_hd__mux2_2
XFILLER_130_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6175_ _9571_/Q _6166_/A _7976_/A _6197_/A vssd1 vssd1 vccd1 vccd1 _6179_/A sky130_fd_sc_hd__a22o_1
X_5126_ _4743_/X _9793_/Q _5121_/X _9220_/X _5124_/X vssd1 vssd1 vccd1 vccd1 _9793_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_84_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5057_ _9809_/Q vssd1 vssd1 vccd1 vccd1 _6316_/C sky130_fd_sc_hd__inv_2
XFILLER_84_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_9865_ _9874_/CLK _9865_/D vssd1 vssd1 vccd1 vccd1 _9865_/Q sky130_fd_sc_hd__dfxtp_1
X_8816_ _8814_/X _8815_/X _8814_/X _8815_/X vssd1 vssd1 vccd1 vccd1 _8816_/X sky130_fd_sc_hd__a2bb2o_1
X_9796_ _9796_/CLK _9796_/D vssd1 vssd1 vccd1 vccd1 _9796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8747_ _8747_/A _8747_/B vssd1 vssd1 vccd1 vccd1 _8797_/A sky130_fd_sc_hd__nand2_1
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5959_ _5959_/A vssd1 vssd1 vccd1 vccd1 _5959_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8678_ _8714_/A _8634_/B _8677_/Y _8634_/Y _8677_/A vssd1 vssd1 vccd1 vccd1 _8678_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_193_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7629_ _7593_/A _7593_/B _7594_/B vssd1 vssd1 vccd1 vccd1 _7629_/X sky130_fd_sc_hd__a21bo_1
XFILLER_193_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7980_ _8980_/X _8002_/B vssd1 vssd1 vccd1 vccd1 _7980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6931_ _6923_/Y _6927_/X _6929_/X _6930_/X vssd1 vssd1 vccd1 vccd1 _6931_/X sky130_fd_sc_hd__o22a_1
XFILLER_207_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9650_ _9650_/CLK _9650_/D vssd1 vssd1 vccd1 vccd1 _9650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6862_ _6862_/A vssd1 vssd1 vccd1 vccd1 _6881_/B sky130_fd_sc_hd__buf_1
XFILLER_179_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8601_ _8387_/X _8404_/X _8387_/X _8404_/X vssd1 vssd1 vccd1 vccd1 _8602_/A sky130_fd_sc_hd__a2bb2o_1
X_9581_ _9833_/CLK _9581_/D vssd1 vssd1 vccd1 vccd1 _9581_/Q sky130_fd_sc_hd__dfxtp_1
X_5813_ _9652_/Q _5557_/X _4900_/X _7083_/B _5809_/X vssd1 vssd1 vccd1 vccd1 _9652_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8532_ _8458_/A _8479_/A _8510_/Y _8508_/A _8531_/Y vssd1 vssd1 vccd1 vccd1 _8532_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_179_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6793_ _6821_/B _6868_/B _6796_/D _6862_/A vssd1 vssd1 vccd1 vccd1 _6795_/A sky130_fd_sc_hd__o22a_1
XFILLER_210_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5744_ _5744_/A vssd1 vssd1 vccd1 vccd1 _5744_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8463_ _8463_/A _8463_/B vssd1 vssd1 vccd1 vccd1 _8486_/A sky130_fd_sc_hd__or2_1
X_5675_ _5515_/X _5671_/X _6804_/C _5662_/X _5674_/X vssd1 vssd1 vccd1 vccd1 _9684_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_175_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8394_ _8394_/A _8394_/B vssd1 vssd1 vccd1 vccd1 _8394_/Y sky130_fd_sc_hd__nor2_1
X_7414_ _7399_/A _7409_/Y _7406_/X _7410_/X vssd1 vssd1 vccd1 vccd1 _7421_/A sky130_fd_sc_hd__o22ai_4
XFILLER_190_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7345_ _7324_/C _7320_/X _7324_/C _7320_/X vssd1 vssd1 vccd1 vccd1 _7346_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_171_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7276_ _7276_/A _7276_/B vssd1 vssd1 vccd1 vccd1 _7276_/X sky130_fd_sc_hd__or2_2
X_9015_ _9783_/Q _9900_/Q _9480_/S vssd1 vssd1 vccd1 vccd1 _9015_/X sky130_fd_sc_hd__mux2_1
X_6227_ _9580_/Q _6168_/A _8015_/A _6241_/A vssd1 vssd1 vccd1 vccd1 _6232_/B sky130_fd_sc_hd__a22o_1
XFILLER_103_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6158_ _9569_/Q vssd1 vssd1 vccd1 vccd1 _7965_/A sky130_fd_sc_hd__inv_2
X_5109_ _9830_/Q vssd1 vssd1 vccd1 vccd1 _5109_/Y sky130_fd_sc_hd__inv_2
X_6089_ _6088_/A _6088_/B _6088_/X vssd1 vssd1 vccd1 vccd1 _6089_/Y sky130_fd_sc_hd__a21boi_1
X_9917_ _9917_/CLK _9917_/D vssd1 vssd1 vccd1 vccd1 _9917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_9848_ _9930_/CLK _9848_/D vssd1 vssd1 vccd1 vccd1 _9848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_9779_ _9898_/CLK _9779_/D vssd1 vssd1 vccd1 vccd1 _9779_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_15_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput52 _9561_/Q vssd1 vssd1 vccd1 vccd1 io_pwm_l sky130_fd_sc_hd__clkbuf_2
XFILLER_122_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput74 _9066_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[28] sky130_fd_sc_hd__clkbuf_2
Xoutput63 _9056_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[18] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput85 _9035_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5460_ _9363_/X _9361_/X _5418_/Y _5483_/A vssd1 vssd1 vccd1 vccd1 _5479_/A sky130_fd_sc_hd__o22a_1
XFILLER_172_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5391_ _5391_/A vssd1 vssd1 vccd1 vccd1 _9720_/D sky130_fd_sc_hd__inv_2
XFILLER_153_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7130_ _7389_/A vssd1 vssd1 vccd1 vccd1 _7385_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_207_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7061_ _7061_/A vssd1 vssd1 vccd1 vccd1 _7076_/A sky130_fd_sc_hd__inv_2
XFILLER_207_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6012_ _9852_/Q _6004_/Y _6009_/A vssd1 vssd1 vccd1 vccd1 _6019_/A sky130_fd_sc_hd__o21ai_1
.ends

